--副程式:OLED
--1. Libraries Declarations and Packages usage
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
--*****************************************************************************
--2. Entity Declarations
entity OLED is 
port(-- input signals
	 clk        : in	std_logic; -- Pin = 149 , 50MHz
	 rst	    : in	std_logic; -- active Low (Internal)
     tft_lcd_p  : in	std_logic; -- 10MHz Pulsed Wave
     start_p    : in	std_logic; -- Tw = 20nS
     rgb_code   : in    integer range 0 to 10; -- Well-defined Color Code
     word_code  : in    integer range 0 to 15; -- Well-defined Color Code
     rgb_color  : in	std_logic_vector(15 downto 0); -- Self Defined Color
     word_color : in	std_logic_vector(15 downto 0); -- Self Defined Color
     data_in    : in	integer range 0 to 82;         -- Digits (BCD Codes)
     row_addr   : in	integer range 0 to 159;        -- 0 ~ 160
     row_range  : in	integer range 1 to 160;
     col_addr   : in	integer range 0 to 127;        -- 0 ~ 127
     col_range  : in	integer range 1 to 128;
     font_sel   : in	integer range 0 to 10;         -- 0 : 32x32 , 1 : 16x16 , 2 : picture
     -- output signals
     bf_out     : out   std_logic; -- 1 : component is busy. ; 0 : Ready
     -- RGB TFT LCD I/O signals
     BL_tft     : out   std_logic; -- active High
     rst_tft    : out   std_logic; -- active Low
     cs         : out   std_logic; -- SPI : active Low , NET , PET
     dc         : out   std_logic; -- SPI : 0 : Command ; 1 : Data
     scl        : out   std_logic; -- SPI : clock
     sda        : out   std_logic  -- SPI : data  line
	);
end OLED;
--*****************************************************************************
--3. Architectures (Body)
architecture beh of OLED is
	-- Global Signals
	signal flag_init  : std_logic_vector( 1 downto 0);
    signal flag_start : std_logic;
    signal code       : std_logic_vector( 7 downto 0);
    signal color_bkgd : std_logic_vector(15 downto 0);
    signal color_word : std_logic_vector(15 downto 0);
    signal color      : std_logic_vector(15 downto 0);
    signal row_y1     : std_logic_vector( 7 downto 0); 
    signal col_x1     : std_logic_vector( 7 downto 0);
    signal row_y2     : std_logic_vector( 7 downto 0);
    signal col_x2     : std_logic_vector( 7 downto 0); 
    signal col_r_8    : integer range 0 to 128;
    signal col_r      : integer range 0 to 128;
    signal row_r      : integer range 0 to 160;
    signal index_t    : integer range 0 to 20480;  
    signal bcd        : integer range 0 to 82;
    signal font_bit   : std_logic;
    signal color_bit  : std_logic;
    ---------------------------------------------------------------------------
    -- Fonts
	-- Dummy Font
    type rom160x128 is array (0 to 2559) of std_logic_vector(7 downto 0);
	constant Font160 : rom160x128 :=( -- 160 x 128 / 8 = 2560 Bytes (rows x cols = H x W)
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00");
	--------------------------------------------------------------------------------
	-- 0~9 A~Z a~z 
    type rom53x32 is array (0 to 82, 0 to 211) of std_logic_vector(7 downto 0); 
	constant Font53 : rom53x32 :=( -- 53 x 32 / 8 = 212 Bytes (rows x cols = H x W)
							   (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 0
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", 
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"07",X"E0",X"00",X"00",X"1F",X"F8",X"00",
								X"00",X"3F",X"FC",X"00",X"00",X"7F",X"FE",X"00",
								X"00",X"FC",X"7F",X"00",X"01",X"F8",X"1F",X"80",
								X"01",X"F0",X"0F",X"80",X"01",X"F0",X"0F",X"80",
								X"03",X"E0",X"07",X"C0",X"03",X"E0",X"0F",X"C0",
								X"03",X"E0",X"1F",X"C0",X"03",X"E0",X"3F",X"C0",
								X"07",X"C0",X"3F",X"C0",X"07",X"C0",X"7B",X"E0",
								X"07",X"C0",X"F3",X"E0",X"07",X"C1",X"E3",X"E0",
								X"07",X"C3",X"C3",X"E0",X"07",X"C7",X"83",X"E0",
								X"07",X"C7",X"83",X"E0",X"07",X"CF",X"03",X"E0",
								X"07",X"DE",X"03",X"E0",X"03",X"FC",X"07",X"C0",
								X"03",X"F8",X"07",X"C0",X"03",X"F0",X"07",X"C0",
								X"03",X"E0",X"07",X"C0",X"01",X"F0",X"0F",X"80",
								X"01",X"F0",X"0F",X"80",X"01",X"F8",X"1F",X"80",
								X"00",X"FC",X"3F",X"00",X"00",X"7F",X"FE",X"00",
								X"00",X"3F",X"FC",X"00",X"00",X"1F",X"F8",X"00",
								X"00",X"07",X"E0",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
							   -------------------------------------------------
							   (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 1
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"01",X"E0",X"00",X"00",X"07",X"E0",X"00",
								X"00",X"1F",X"E0",X"00",X"00",X"7F",X"E0",X"00",
								X"01",X"FF",X"E0",X"00",X"01",X"FF",X"E0",X"00",
								X"00",X"F3",X"E0",X"00",X"00",X"83",X"E0",X"00",
								X"00",X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",
								X"00",X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",
								X"00",X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",
								X"00",X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",
								X"00",X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",
								X"00",X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",
								X"00",X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",
								X"00",X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",
								X"00",X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",
								X"00",X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",
								X"00",X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",
								X"00",X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
							   -------------------------------------------------
							   (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 2
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"07",X"F0",X"00",X"00",X"3F",X"FC",X"00",
								X"00",X"7F",X"FE",X"00",X"01",X"FF",X"FF",X"00",
								X"01",X"FE",X"7F",X"80",X"03",X"F0",X"0F",X"80",
								X"03",X"E0",X"0F",X"C0",X"01",X"C0",X"07",X"C0",
								X"00",X"C0",X"07",X"C0",X"00",X"00",X"07",X"C0",
								X"00",X"00",X"07",X"C0",X"00",X"00",X"07",X"C0",
								X"00",X"00",X"0F",X"80",X"00",X"00",X"0F",X"80",
								X"00",X"00",X"1F",X"80",X"00",X"00",X"1F",X"00",
								X"00",X"00",X"3E",X"00",X"00",X"00",X"7E",X"00",
								X"00",X"00",X"FC",X"00",X"00",X"01",X"F8",X"00",
								X"00",X"03",X"F0",X"00",X"00",X"07",X"E0",X"00",
								X"00",X"0F",X"C0",X"00",X"00",X"1F",X"80",X"00",
								X"00",X"3F",X"00",X"00",X"00",X"7E",X"00",X"00",
								X"00",X"FC",X"00",X"00",X"01",X"F8",X"00",X"40",
								X"03",X"FF",X"FF",X"C0",X"03",X"FF",X"FF",X"C0",
								X"03",X"FF",X"FF",X"C0",X"03",X"FF",X"FF",X"C0",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
							   -------------------------------------------------
							   (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 3
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"0F",X"E0",X"00",X"00",X"7F",X"F8",X"00",
								X"00",X"FF",X"FC",X"00",X"01",X"FF",X"FE",X"00",
								X"01",X"F8",X"7F",X"00",X"00",X"E0",X"1F",X"00",
								X"00",X"40",X"1F",X"80",X"00",X"00",X"0F",X"80",
								X"00",X"00",X"0F",X"80",X"00",X"00",X"0F",X"80",
								X"00",X"00",X"1F",X"00",X"00",X"00",X"1F",X"00",
								X"00",X"00",X"3F",X"00",X"00",X"00",X"FE",X"00",
								X"00",X"0F",X"FC",X"00",X"00",X"0F",X"F0",X"00",
								X"00",X"0F",X"FC",X"00",X"00",X"0F",X"FE",X"00",
								X"00",X"00",X"7F",X"00",X"00",X"00",X"1F",X"80",
								X"00",X"00",X"0F",X"80",X"00",X"00",X"0F",X"80",
								X"00",X"00",X"0F",X"C0",X"00",X"00",X"07",X"C0",
								X"00",X"00",X"0F",X"C0",X"00",X"80",X"0F",X"C0",
								X"00",X"C0",X"0F",X"80",X"01",X"E0",X"1F",X"80",
								X"03",X"F8",X"7F",X"00",X"03",X"FF",X"FF",X"00",
								X"01",X"FF",X"FE",X"00",X"00",X"7F",X"F8",X"00",
								X"00",X"1F",X"E0",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
							   -------------------------------------------------
							   (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 4
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 4
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"1E",X"00",X"00",X"00",X"3E",X"00",
								X"00",X"00",X"3E",X"00",X"00",X"00",X"7E",X"00",
								X"00",X"00",X"FE",X"00",X"00",X"00",X"FE",X"00",
								X"00",X"01",X"FE",X"00",X"00",X"03",X"FE",X"00",
								X"00",X"03",X"FE",X"00",X"00",X"07",X"FE",X"00",
								X"00",X"0F",X"BE",X"00",X"00",X"1F",X"3E",X"00",
								X"00",X"1E",X"3E",X"00",X"00",X"3E",X"3E",X"00",
								X"00",X"7C",X"3E",X"00",X"00",X"78",X"3E",X"00",
								X"00",X"F8",X"3E",X"00",X"01",X"F0",X"3E",X"00",
								X"01",X"E0",X"3E",X"00",X"03",X"E0",X"3E",X"00",
								X"07",X"FF",X"FF",X"F0",X"07",X"FF",X"FF",X"F0",
								X"07",X"FF",X"FF",X"F0",X"07",X"FF",X"FF",X"F0",
								X"00",X"00",X"3E",X"00",X"00",X"00",X"3E",X"00",
								X"00",X"00",X"3E",X"00",X"00",X"00",X"3E",X"00",
								X"00",X"00",X"3E",X"00",X"00",X"00",X"3E",X"00",
								X"00",X"00",X"3E",X"00",X"00",X"00",X"3E",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
							   -------------------------------------------------
							   (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 5
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 5
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"FF",X"FF",X"80",X"00",X"FF",X"FF",X"80",
								X"00",X"FF",X"FF",X"80",X"00",X"FF",X"FF",X"80",
								X"00",X"F8",X"00",X"00",X"00",X"F8",X"00",X"00",
								X"00",X"F8",X"00",X"00",X"00",X"F0",X"00",X"00",
								X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",
								X"00",X"F0",X"00",X"00",X"00",X"F3",X"F0",X"00",
								X"01",X"FF",X"FC",X"00",X"01",X"FF",X"FF",X"00",
								X"01",X"FF",X"FF",X"00",X"01",X"FC",X"3F",X"80",
								X"01",X"F0",X"0F",X"C0",X"00",X"60",X"0F",X"C0",
								X"00",X"00",X"07",X"C0",X"00",X"00",X"07",X"C0",
								X"00",X"00",X"03",X"E0",X"00",X"00",X"03",X"E0",
								X"00",X"00",X"03",X"E0",X"00",X"00",X"03",X"E0",
								X"00",X"00",X"07",X"C0",X"00",X"40",X"07",X"C0",
								X"00",X"E0",X"0F",X"C0",X"03",X"F0",X"1F",X"80",
								X"03",X"FC",X"3F",X"80",X"01",X"FF",X"FF",X"00",
								X"00",X"FF",X"FE",X"00",X"00",X"3F",X"FC",X"00",
								X"00",X"0F",X"E0",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
							   -------------------------------------------------
							   (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 6
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 6
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"01",X"F8",X"00",X"00",X"07",X"FF",X"00",
								X"00",X"1F",X"FF",X"80",X"00",X"3F",X"FF",X"80",
								X"00",X"7F",X"8F",X"00",X"00",X"7E",X"03",X"00",
								X"00",X"FC",X"02",X"00",X"00",X"F8",X"00",X"00",
								X"01",X"F0",X"00",X"00",X"01",X"F0",X"00",X"00",
								X"01",X"F0",X"00",X"00",X"01",X"E0",X"00",X"00",
								X"03",X"E1",X"F0",X"00",X"03",X"E7",X"FC",X"00",
								X"03",X"EF",X"FF",X"00",X"03",X"FF",X"FF",X"00",
								X"03",X"FE",X"3F",X"80",X"03",X"F8",X"0F",X"C0",
								X"03",X"F0",X"07",X"C0",X"03",X"E0",X"07",X"C0",
								X"03",X"E0",X"07",X"C0",X"03",X"E0",X"03",X"C0",
								X"03",X"E0",X"03",X"C0",X"01",X"E0",X"07",X"C0",
								X"01",X"F0",X"07",X"C0",X"01",X"F0",X"07",X"C0",
								X"01",X"F8",X"0F",X"C0",X"00",X"FC",X"0F",X"80",
								X"00",X"FE",X"3F",X"80",X"00",X"7F",X"FF",X"00",
								X"00",X"3F",X"FE",X"00",X"00",X"1F",X"FC",X"00",
								X"00",X"07",X"F0",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
							   -------------------------------------------------
							   (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 7
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 7
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"01",X"FF",X"FF",X"C0",X"01",X"FF",X"FF",X"C0",
								X"01",X"FF",X"FF",X"C0",X"01",X"FF",X"FF",X"C0",
								X"01",X"FF",X"FF",X"80",X"00",X"00",X"1F",X"80",
								X"00",X"00",X"1F",X"00",X"00",X"00",X"1F",X"00",
								X"00",X"00",X"3F",X"00",X"00",X"00",X"3E",X"00",
								X"00",X"00",X"3E",X"00",X"00",X"00",X"7C",X"00",
								X"00",X"00",X"7C",X"00",X"00",X"00",X"FC",X"00",
								X"00",X"00",X"F8",X"00",X"00",X"00",X"F8",X"00",
								X"00",X"01",X"F0",X"00",X"00",X"01",X"F0",X"00",
								X"00",X"01",X"F0",X"00",X"00",X"03",X"E0",X"00",
								X"00",X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",
								X"00",X"07",X"C0",X"00",X"00",X"07",X"C0",X"00",
								X"00",X"0F",X"C0",X"00",X"00",X"0F",X"80",X"00",
								X"00",X"0F",X"80",X"00",X"00",X"1F",X"80",X"00",
								X"00",X"1F",X"00",X"00",X"00",X"1F",X"00",X"00",
								X"00",X"3F",X"00",X"00",X"00",X"3F",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
							   -------------------------------------------------
							   (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 8
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 8
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"07",X"F0",X"00",X"00",X"1F",X"FC",X"00",
								X"00",X"7F",X"FE",X"00",X"00",X"7F",X"FF",X"00",
								X"00",X"FC",X"3F",X"80",X"01",X"F8",X"1F",X"80",
								X"01",X"F0",X"0F",X"80",X"01",X"F0",X"0F",X"80",
								X"01",X"F0",X"07",X"80",X"01",X"F0",X"0F",X"80",
								X"01",X"F8",X"0F",X"80",X"00",X"F8",X"1F",X"80",
								X"00",X"FE",X"1F",X"00",X"00",X"7F",X"3E",X"00",
								X"00",X"3F",X"FC",X"00",X"00",X"0F",X"F8",X"00",
								X"00",X"3F",X"FC",X"00",X"00",X"7F",X"FF",X"00",
								X"00",X"F8",X"3F",X"80",X"01",X"F0",X"1F",X"80",
								X"03",X"F0",X"0F",X"C0",X"03",X"E0",X"07",X"C0",
								X"03",X"E0",X"07",X"C0",X"03",X"E0",X"07",X"C0",
								X"03",X"E0",X"07",X"C0",X"03",X"E0",X"07",X"C0",
								X"03",X"F0",X"07",X"C0",X"03",X"F0",X"0F",X"C0",
								X"01",X"FE",X"7F",X"80",X"01",X"FF",X"FF",X"80",
								X"00",X"FF",X"FF",X"00",X"00",X"3F",X"FC",X"00",
								X"00",X"0F",X"F0",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
							   -------------------------------------------------
							   (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 9
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 9
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"07",X"E0",X"00",X"00",X"1F",X"F8",X"00",
								X"00",X"7F",X"FC",X"00",X"00",X"FF",X"FE",X"00",
								X"00",X"FC",X"3F",X"00",X"01",X"F8",X"1F",X"00",
								X"01",X"F0",X"0F",X"80",X"03",X"E0",X"0F",X"80",
								X"03",X"E0",X"07",X"80",X"03",X"E0",X"07",X"C0",
								X"03",X"E0",X"07",X"C0",X"03",X"E0",X"07",X"C0",
								X"03",X"E0",X"07",X"C0",X"03",X"E0",X"07",X"C0",
								X"03",X"F0",X"07",X"C0",X"01",X"F0",X"0F",X"C0",
								X"01",X"FC",X"3F",X"C0",X"00",X"FF",X"FF",X"C0",
								X"00",X"7F",X"FF",X"C0",X"00",X"3F",X"FF",X"C0",
								X"00",X"0F",X"E7",X"C0",X"00",X"00",X"07",X"C0",
								X"00",X"00",X"07",X"80",X"00",X"00",X"0F",X"80",
								X"00",X"00",X"0F",X"80",X"00",X"00",X"1F",X"00",
								X"00",X"40",X"1F",X"00",X"00",X"C0",X"3F",X"00",
								X"01",X"F0",X"FE",X"00",X"01",X"FF",X"FC",X"00",
								X"01",X"FF",X"F8",X"00",X"00",X"FF",X"F0",X"00",
								X"00",X"1F",X"C0",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
							   -------------------------------------------------
							   (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- A
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 10
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"01",X"80",X"00",X"00",X"03",X"C0",X"00",
								X"00",X"03",X"C0",X"00",X"00",X"03",X"C0",X"00",
								X"00",X"07",X"E0",X"00",X"00",X"07",X"E0",X"00",
								X"00",X"07",X"E0",X"00",X"00",X"0F",X"F0",X"00",
								X"00",X"0F",X"F0",X"00",X"00",X"0F",X"F0",X"00",
								X"00",X"1F",X"F8",X"00",X"00",X"1E",X"78",X"00",
								X"00",X"1E",X"78",X"00",X"00",X"3E",X"7C",X"00",
								X"00",X"3C",X"3C",X"00",X"00",X"3C",X"3E",X"00",
								X"00",X"7C",X"3E",X"00",X"00",X"7C",X"3E",X"00",
								X"00",X"F8",X"1F",X"00",X"00",X"F8",X"1F",X"00",
								X"00",X"FF",X"FF",X"00",X"01",X"FF",X"FF",X"80",
								X"01",X"FF",X"FF",X"80",X"01",X"FF",X"FF",X"80",
								X"03",X"E0",X"07",X"C0",X"03",X"E0",X"07",X"C0",
								X"03",X"E0",X"07",X"C0",X"07",X"C0",X"03",X"E0",
								X"07",X"C0",X"03",X"E0",X"07",X"C0",X"03",X"E0",
								X"0F",X"80",X"01",X"F0",X"0F",X"80",X"01",X"F0",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
							    -------------------------------------------------
							   (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- B
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 11
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"07",X"FF",X"F0",X"00",X"07",X"FF",X"FC",X"00",
								X"07",X"FF",X"FF",X"00",X"07",X"FF",X"FF",X"80",
								X"07",X"C0",X"7F",X"80",X"07",X"C0",X"0F",X"C0",
								X"07",X"C0",X"0F",X"C0",X"07",X"C0",X"07",X"C0",
								X"07",X"C0",X"07",X"C0",X"07",X"C0",X"07",X"C0",
								X"07",X"C0",X"0F",X"C0",X"07",X"C0",X"0F",X"80",
								X"07",X"C0",X"7F",X"00",X"07",X"FF",X"FF",X"00",
								X"07",X"FF",X"FC",X"00",X"07",X"FF",X"FE",X"00",
								X"07",X"FF",X"FF",X"00",X"07",X"C0",X"3F",X"80",
								X"07",X"C0",X"0F",X"C0",X"07",X"C0",X"07",X"C0",
								X"07",X"C0",X"03",X"E0",X"07",X"C0",X"03",X"E0",
								X"07",X"C0",X"03",X"E0",X"07",X"C0",X"03",X"E0",
								X"07",X"C0",X"03",X"E0",X"07",X"C0",X"07",X"E0",
								X"07",X"C0",X"0F",X"E0",X"07",X"C0",X"7F",X"C0",
								X"07",X"FF",X"FF",X"80",X"07",X"FF",X"FF",X"00",
								X"07",X"FF",X"FE",X"00",X"07",X"FF",X"F0",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
							    -------------------------------------------------
							   (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- C
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 12
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"03",X"F8",X"00",X"00",X"0F",X"FF",X"00",
								X"00",X"3F",X"FF",X"80",X"00",X"7F",X"FF",X"C0",
								X"00",X"FF",X"0F",X"E0",X"01",X"FC",X"03",X"E0",
								X"01",X"F8",X"01",X"F0",X"03",X"F0",X"01",X"C0",
								X"03",X"E0",X"00",X"80",X"03",X"E0",X"00",X"00",
								X"07",X"E0",X"00",X"00",X"07",X"C0",X"00",X"00",
								X"07",X"C0",X"00",X"00",X"07",X"C0",X"00",X"00",
								X"07",X"C0",X"00",X"00",X"07",X"C0",X"00",X"00",
								X"07",X"C0",X"00",X"00",X"07",X"C0",X"00",X"00",
								X"07",X"C0",X"00",X"00",X"07",X"C0",X"00",X"00",
								X"07",X"C0",X"00",X"00",X"07",X"C0",X"00",X"00",
								X"07",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"F0",X"00",X"00",X"03",X"F0",X"01",X"00",
								X"01",X"F8",X"01",X"C0",X"01",X"FC",X"03",X"E0",
								X"00",X"FF",X"1F",X"E0",X"00",X"7F",X"FF",X"C0",
								X"00",X"3F",X"FF",X"80",X"00",X"0F",X"FF",X"00",
								X"00",X"03",X"F8",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
							    -------------------------------------------------
							   (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- D
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 13
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"07",X"FF",X"C0",X"00",X"07",X"FF",X"F8",X"00",
								X"07",X"FF",X"FC",X"00",X"07",X"FF",X"FE",X"00",
								X"07",X"C0",X"FF",X"00",X"07",X"C0",X"3F",X"80",
								X"07",X"C0",X"0F",X"80",X"07",X"C0",X"0F",X"C0",
								X"07",X"C0",X"07",X"C0",X"07",X"C0",X"07",X"C0",
								X"07",X"C0",X"03",X"E0",X"07",X"C0",X"03",X"E0",
								X"07",X"C0",X"03",X"E0",X"07",X"C0",X"03",X"E0",
								X"07",X"C0",X"03",X"E0",X"07",X"C0",X"03",X"E0",
								X"07",X"C0",X"03",X"E0",X"07",X"C0",X"03",X"E0",
								X"07",X"C0",X"03",X"E0",X"07",X"C0",X"03",X"E0",
								X"07",X"C0",X"03",X"E0",X"07",X"C0",X"03",X"E0",
								X"07",X"C0",X"07",X"E0",X"07",X"C0",X"07",X"C0",
								X"07",X"C0",X"0F",X"C0",X"07",X"C0",X"0F",X"80",
								X"07",X"C0",X"3F",X"80",X"07",X"C0",X"FF",X"00",
								X"07",X"FF",X"FE",X"00",X"07",X"FF",X"FC",X"00",
								X"07",X"FF",X"F0",X"00",X"07",X"FF",X"80",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- E
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 14
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"03",X"FF",X"FF",X"C0",X"03",X"FF",X"FF",X"C0",
								X"03",X"FF",X"FF",X"C0",X"03",X"FF",X"FF",X"C0",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"FF",X"FF",X"00",
								X"03",X"FF",X"FF",X"00",X"03",X"FF",X"FF",X"00",
								X"03",X"FF",X"FF",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"FF",X"FF",X"C0",X"03",X"FF",X"FF",X"C0",
								X"03",X"FF",X"FF",X"C0",X"03",X"FF",X"FF",X"C0",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- F
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 15
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"01",X"FF",X"FF",X"C0",X"01",X"FF",X"FF",X"C0",
								X"01",X"FF",X"FF",X"C0",X"01",X"FF",X"FF",X"C0",
								X"01",X"E0",X"00",X"00",X"01",X"E0",X"00",X"00",
								X"01",X"E0",X"00",X"00",X"01",X"E0",X"00",X"00",
								X"01",X"E0",X"00",X"00",X"01",X"E0",X"00",X"00",
								X"01",X"E0",X"00",X"00",X"01",X"E0",X"00",X"00",
								X"01",X"E0",X"00",X"00",X"01",X"FF",X"FE",X"00",
								X"01",X"FF",X"FE",X"00",X"01",X"FF",X"FE",X"00",
								X"01",X"FF",X"FE",X"00",X"01",X"E0",X"00",X"00",
								X"01",X"E0",X"00",X"00",X"01",X"E0",X"00",X"00",
								X"01",X"E0",X"00",X"00",X"01",X"E0",X"00",X"00",
								X"01",X"E0",X"00",X"00",X"01",X"E0",X"00",X"00",
								X"01",X"E0",X"00",X"00",X"01",X"E0",X"00",X"00",
								X"01",X"E0",X"00",X"00",X"01",X"E0",X"00",X"00",
								X"01",X"E0",X"00",X"00",X"01",X"E0",X"00",X"00",
								X"01",X"E0",X"00",X"00",X"01",X"E0",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- G
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 16
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"03",X"F8",X"00",X"00",X"1F",X"FE",X"00",
								X"00",X"3F",X"FF",X"80",X"00",X"7F",X"FF",X"C0",
								X"00",X"FF",X"1F",X"E0",X"01",X"F8",X"07",X"E0",
								X"01",X"F0",X"03",X"C0",X"03",X"F0",X"01",X"80",
								X"03",X"E0",X"01",X"00",X"07",X"E0",X"00",X"00",
								X"07",X"C0",X"00",X"00",X"07",X"C0",X"00",X"00",
								X"07",X"C0",X"00",X"00",X"07",X"C0",X"00",X"00",
								X"07",X"C0",X"00",X"00",X"0F",X"C0",X"00",X"00",
								X"07",X"C0",X"00",X"00",X"07",X"C0",X"7F",X"E0",
								X"07",X"C0",X"7F",X"E0",X"07",X"C0",X"7F",X"E0",
								X"07",X"C0",X"7F",X"E0",X"07",X"C0",X"01",X"E0",
								X"07",X"C0",X"01",X"E0",X"07",X"E0",X"01",X"E0",
								X"03",X"E0",X"01",X"E0",X"03",X"F0",X"01",X"E0",
								X"01",X"F0",X"01",X"E0",X"01",X"FC",X"03",X"E0",
								X"00",X"FF",X"1F",X"E0",X"00",X"7F",X"FF",X"E0",
								X"00",X"3F",X"FF",X"C0",X"00",X"1F",X"FF",X"00",
								X"00",X"03",X"F8",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- H
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 17
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"07",X"E0",X"07",X"E0",X"07",X"C0",X"07",X"E0",
								X"07",X"C0",X"07",X"E0",X"07",X"C0",X"07",X"E0",
								X"07",X"C0",X"07",X"E0",X"07",X"C0",X"07",X"E0",
								X"07",X"C0",X"07",X"E0",X"07",X"C0",X"07",X"E0",
								X"07",X"C0",X"07",X"E0",X"07",X"C0",X"07",X"E0",
								X"07",X"C0",X"07",X"E0",X"07",X"C0",X"07",X"E0",
								X"07",X"C0",X"07",X"E0",X"07",X"FF",X"FF",X"E0",
								X"07",X"FF",X"FF",X"E0",X"07",X"FF",X"FF",X"E0",
								X"07",X"FF",X"FF",X"E0",X"07",X"C0",X"07",X"E0",
								X"07",X"C0",X"07",X"E0",X"07",X"C0",X"07",X"E0",
								X"07",X"C0",X"07",X"E0",X"07",X"C0",X"07",X"E0",
								X"07",X"C0",X"07",X"E0",X"07",X"C0",X"07",X"E0",
								X"07",X"C0",X"07",X"E0",X"07",X"C0",X"07",X"E0",
								X"07",X"C0",X"07",X"E0",X"07",X"C0",X"07",X"E0",
								X"07",X"C0",X"07",X"E0",X"07",X"C0",X"07",X"E0",
								X"07",X"C0",X"07",X"E0",X"07",X"C0",X"07",X"E0",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- I
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 18
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"01",X"FF",X"FF",X"00",X"01",X"FF",X"FF",X"00",
								X"01",X"FF",X"FF",X"00",X"01",X"FF",X"FF",X"00",
								X"00",X"07",X"C0",X"00",X"00",X"07",X"C0",X"00",
								X"00",X"07",X"C0",X"00",X"00",X"07",X"C0",X"00",
								X"00",X"07",X"C0",X"00",X"00",X"07",X"C0",X"00",
								X"00",X"07",X"C0",X"00",X"00",X"07",X"C0",X"00",
								X"00",X"07",X"C0",X"00",X"00",X"07",X"C0",X"00",
								X"00",X"07",X"C0",X"00",X"00",X"07",X"C0",X"00",
								X"00",X"07",X"C0",X"00",X"00",X"07",X"C0",X"00",
								X"00",X"07",X"C0",X"00",X"00",X"07",X"C0",X"00",
								X"00",X"07",X"C0",X"00",X"00",X"07",X"C0",X"00",
								X"00",X"07",X"C0",X"00",X"00",X"07",X"C0",X"00",
								X"00",X"07",X"C0",X"00",X"00",X"07",X"C0",X"00",
								X"00",X"07",X"C0",X"00",X"00",X"07",X"C0",X"00",
								X"01",X"FF",X"FF",X"80",X"01",X"FF",X"FF",X"80",
								X"01",X"FF",X"FF",X"80",X"01",X"FF",X"FF",X"80",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- J
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 19
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"1F",X"FF",X"E0",X"00",X"1F",X"FF",X"E0",
								X"00",X"1F",X"FF",X"E0",X"00",X"1F",X"FF",X"E0",
								X"00",X"00",X"7C",X"00",X"00",X"00",X"7C",X"00",
								X"00",X"00",X"7C",X"00",X"00",X"00",X"7C",X"00",
								X"00",X"00",X"7C",X"00",X"00",X"00",X"7C",X"00",
								X"00",X"00",X"7C",X"00",X"00",X"00",X"7C",X"00",
								X"00",X"00",X"7C",X"00",X"00",X"00",X"7C",X"00",
								X"00",X"00",X"7C",X"00",X"00",X"00",X"7C",X"00",
								X"00",X"00",X"7C",X"00",X"00",X"00",X"7C",X"00",
								X"00",X"00",X"7C",X"00",X"00",X"00",X"7C",X"00",
								X"00",X"00",X"7C",X"00",X"00",X"00",X"7C",X"00",
								X"00",X"00",X"7C",X"00",X"00",X"00",X"7C",X"00",
								X"00",X"00",X"7C",X"00",X"00",X"00",X"7C",X"00",
								X"01",X"80",X"FC",X"00",X"03",X"C1",X"F8",X"00",
								X"03",X"FF",X"F8",X"00",X"07",X"FF",X"F0",X"00",
								X"03",X"FF",X"E0",X"00",X"01",X"FF",X"C0",X"00",
								X"00",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- K
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 20
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"07",X"E0",X"07",X"E0",
								X"07",X"C0",X"0F",X"C0",X"07",X"C0",X"0F",X"80",
								X"07",X"C0",X"1F",X"80",X"07",X"C0",X"3F",X"00",
								X"07",X"C0",X"7E",X"00",X"07",X"C0",X"FC",X"00",
								X"07",X"C1",X"F8",X"00",X"07",X"C3",X"F0",X"00",
								X"07",X"C3",X"F0",X"00",X"07",X"C7",X"E0",X"00",
								X"07",X"CF",X"C0",X"00",X"07",X"DF",X"80",X"00",
								X"07",X"FF",X"00",X"00",X"07",X"FF",X"80",X"00",
								X"07",X"FF",X"80",X"00",X"07",X"FF",X"C0",X"00",
								X"07",X"F7",X"E0",X"00",X"07",X"E7",X"E0",X"00",
								X"07",X"C3",X"F0",X"00",X"07",X"C1",X"F8",X"00",
								X"07",X"C1",X"F8",X"00",X"07",X"C0",X"FC",X"00",
								X"07",X"C0",X"7E",X"00",X"07",X"C0",X"7E",X"00",
								X"07",X"C0",X"3F",X"00",X"07",X"C0",X"1F",X"80",
								X"07",X"C0",X"1F",X"80",X"07",X"C0",X"0F",X"C0",
								X"07",X"C0",X"0F",X"E0",X"07",X"C0",X"07",X"E0",
								X"07",X"C0",X"03",X"F0",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- L
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 21
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"03",X"F0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"FF",X"FF",X"C0",X"03",X"FF",X"FF",X"C0",
								X"03",X"FF",X"FF",X"C0",X"03",X"FF",X"FF",X"C0",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- M
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 22
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"07",X"80",X"01",X"E0",
								X"07",X"C0",X"03",X"E0",X"07",X"C0",X"03",X"E0",
								X"07",X"E0",X"07",X"E0",X"07",X"E0",X"07",X"E0",
								X"07",X"F0",X"0F",X"E0",X"07",X"F0",X"0F",X"E0",
								X"07",X"F8",X"0F",X"E0",X"07",X"F8",X"1F",X"E0",
								X"07",X"FC",X"1F",X"E0",X"07",X"BC",X"3D",X"E0",
								X"07",X"BC",X"3D",X"E0",X"07",X"9E",X"79",X"E0",
								X"07",X"9E",X"79",X"E0",X"07",X"8F",X"F1",X"E0",
								X"07",X"8F",X"F1",X"E0",X"07",X"87",X"E1",X"E0",
								X"07",X"87",X"E1",X"E0",X"07",X"87",X"C1",X"E0",
								X"07",X"83",X"C1",X"E0",X"07",X"83",X"81",X"E0",
								X"07",X"80",X"01",X"E0",X"07",X"80",X"01",X"E0",
								X"07",X"80",X"01",X"E0",X"07",X"80",X"01",X"E0",
								X"07",X"80",X"01",X"E0",X"07",X"80",X"01",X"E0",
								X"07",X"80",X"01",X"E0",X"07",X"80",X"01",X"E0",
								X"07",X"80",X"01",X"E0",X"07",X"80",X"01",X"E0",
								X"07",X"80",X"01",X"E0",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- N
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 23
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"07",X"E0",X"03",X"E0",X"07",X"E0",X"03",X"E0",
								X"07",X"F0",X"03",X"E0",X"07",X"F0",X"03",X"E0",
								X"07",X"F8",X"03",X"E0",X"07",X"F8",X"03",X"E0",
								X"07",X"FC",X"03",X"E0",X"07",X"FC",X"03",X"E0",
								X"07",X"FE",X"03",X"E0",X"07",X"FF",X"03",X"E0",
								X"07",X"DF",X"03",X"E0",X"07",X"DF",X"83",X"E0",
								X"07",X"CF",X"83",X"E0",X"07",X"CF",X"C3",X"E0",
								X"07",X"C7",X"C3",X"E0",X"07",X"C7",X"E3",X"E0",
								X"07",X"C3",X"E3",X"E0",X"07",X"C3",X"F3",X"E0",
								X"07",X"C1",X"F3",X"E0",X"07",X"C0",X"FB",X"E0",
								X"07",X"C0",X"FF",X"E0",X"07",X"C0",X"7F",X"E0",
								X"07",X"C0",X"7F",X"E0",X"07",X"C0",X"3F",X"E0",
								X"07",X"C0",X"3F",X"E0",X"07",X"C0",X"1F",X"E0",
								X"07",X"C0",X"1F",X"E0",X"07",X"C0",X"0F",X"E0",
								X"07",X"C0",X"0F",X"E0",X"07",X"C0",X"07",X"E0",
								X"07",X"C0",X"07",X"E0",X"07",X"C0",X"03",X"E0",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- O
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 24
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"0F",X"F0",X"00",X"00",X"3F",X"FC",X"00",
								X"00",X"7F",X"FE",X"00",X"00",X"FF",X"FF",X"00",
								X"01",X"FE",X"3F",X"80",X"03",X"F8",X"1F",X"C0",
								X"03",X"F0",X"0F",X"C0",X"03",X"E0",X"07",X"E0",
								X"07",X"E0",X"03",X"E0",X"07",X"C0",X"03",X"E0",
								X"07",X"C0",X"03",X"E0",X"0F",X"C0",X"03",X"F0",
								X"0F",X"C0",X"01",X"F0",X"0F",X"80",X"01",X"F0",
								X"0F",X"80",X"01",X"F0",X"0F",X"80",X"01",X"F0",
								X"0F",X"80",X"01",X"F0",X"0F",X"80",X"01",X"F0",
								X"0F",X"80",X"01",X"F0",X"0F",X"80",X"01",X"F0",
								X"0F",X"C0",X"01",X"F0",X"0F",X"C0",X"03",X"F0",
								X"07",X"C0",X"03",X"E0",X"07",X"C0",X"03",X"E0",
								X"07",X"C0",X"03",X"E0",X"07",X"E0",X"07",X"E0",
								X"03",X"F0",X"0F",X"C0",X"03",X"F8",X"0F",X"C0",
								X"01",X"FC",X"3F",X"80",X"00",X"FF",X"FF",X"00",
								X"00",X"7F",X"FE",X"00",X"00",X"3F",X"FC",X"00",
								X"00",X"0F",X"F0",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- P
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 25
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"03",X"FF",X"F8",X"00",X"03",X"FF",X"FE",X"00",
								X"03",X"FF",X"FF",X"00",X"03",X"FF",X"FF",X"80",
								X"03",X"FF",X"FF",X"C0",X"03",X"E0",X"0F",X"E0",
								X"03",X"E0",X"07",X"E0",X"03",X"E0",X"03",X"E0",
								X"03",X"E0",X"03",X"E0",X"03",X"E0",X"03",X"E0",
								X"03",X"E0",X"03",X"E0",X"03",X"E0",X"07",X"E0",
								X"03",X"E0",X"0F",X"E0",X"03",X"E0",X"3F",X"C0",
								X"03",X"FF",X"FF",X"C0",X"03",X"FF",X"FF",X"80",
								X"03",X"FF",X"FE",X"00",X"03",X"FF",X"F8",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- Q
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 26
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"07",X"E0",X"00",X"00",X"1F",X"FC",X"00",
								X"00",X"7F",X"FE",X"00",X"00",X"FF",X"FF",X"00",
								X"01",X"FC",X"3F",X"80",X"01",X"F8",X"1F",X"C0",
								X"03",X"F0",X"0F",X"C0",X"03",X"E0",X"07",X"C0",
								X"07",X"E0",X"03",X"E0",X"07",X"C0",X"03",X"E0",
								X"07",X"C0",X"03",X"E0",X"07",X"C0",X"03",X"F0",
								X"0F",X"80",X"01",X"F0",X"0F",X"80",X"01",X"F0",
								X"0F",X"80",X"01",X"F0",X"0F",X"80",X"01",X"F0",
								X"0F",X"80",X"01",X"F0",X"0F",X"80",X"01",X"F0",
								X"0F",X"80",X"01",X"F0",X"0F",X"80",X"01",X"F0",
								X"0F",X"80",X"01",X"F0",X"07",X"C0",X"01",X"F0",
								X"07",X"C0",X"03",X"E0",X"07",X"C0",X"03",X"E0",
								X"07",X"E0",X"03",X"E0",X"03",X"E0",X"07",X"E0",
								X"03",X"F0",X"07",X"C0",X"01",X"F8",X"0F",X"C0",
								X"01",X"FC",X"3F",X"80",X"00",X"FF",X"FF",X"00",
								X"00",X"7F",X"FE",X"00",X"00",X"3F",X"FC",X"00",
								X"00",X"0F",X"F0",X"00",X"00",X"03",X"E0",X"00",
								X"00",X"03",X"E0",X"00",X"00",X"03",X"F0",X"00",
								X"00",X"03",X"FF",X"C0",X"00",X"01",X"FF",X"C0",
								X"00",X"00",X"FF",X"C0",X"00",X"00",X"3F",X"C0",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- R
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 27
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"07",X"FF",X"F0",X"00",X"07",X"FF",X"FE",X"00",
								X"07",X"FF",X"FF",X"00",X"07",X"FF",X"FF",X"80",
								X"07",X"FF",X"FF",X"C0",X"07",X"E0",X"0F",X"C0",
								X"07",X"E0",X"07",X"C0",X"07",X"E0",X"07",X"E0",
								X"07",X"E0",X"07",X"E0",X"07",X"E0",X"07",X"E0",
								X"07",X"E0",X"07",X"E0",X"07",X"E0",X"07",X"C0",
								X"07",X"E0",X"0F",X"C0",X"07",X"E0",X"7F",X"C0",
								X"07",X"FF",X"FF",X"80",X"07",X"FF",X"FF",X"00",
								X"07",X"FF",X"FE",X"00",X"07",X"FF",X"F8",X"00",
								X"07",X"E0",X"F8",X"00",X"07",X"E0",X"F8",X"00",
								X"07",X"E0",X"7C",X"00",X"07",X"E0",X"7C",X"00",
								X"07",X"E0",X"3E",X"00",X"07",X"E0",X"3E",X"00",
								X"07",X"E0",X"1F",X"00",X"07",X"E0",X"1F",X"00",
								X"07",X"E0",X"0F",X"80",X"07",X"E0",X"0F",X"80",
								X"07",X"E0",X"0F",X"C0",X"07",X"E0",X"07",X"C0",
								X"07",X"E0",X"07",X"E0",X"07",X"E0",X"03",X"E0",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- S
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 28
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"07",X"F0",X"00",X"00",X"3F",X"FE",X"00",
								X"00",X"7F",X"FF",X"00",X"00",X"FF",X"FF",X"80",
								X"01",X"FC",X"3F",X"C0",X"01",X"F8",X"07",X"80",
								X"03",X"F0",X"03",X"00",X"03",X"E0",X"02",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"F0",X"00",X"00",
								X"01",X"F0",X"00",X"00",X"01",X"F8",X"00",X"00",
								X"01",X"FE",X"00",X"00",X"00",X"FF",X"80",X"00",
								X"00",X"7F",X"E0",X"00",X"00",X"3F",X"F8",X"00",
								X"00",X"0F",X"FE",X"00",X"00",X"03",X"FF",X"00",
								X"00",X"00",X"FF",X"80",X"00",X"00",X"3F",X"C0",
								X"00",X"00",X"0F",X"C0",X"00",X"00",X"07",X"E0",
								X"00",X"00",X"03",X"E0",X"00",X"00",X"03",X"E0",
								X"00",X"00",X"03",X"E0",X"01",X"80",X"03",X"E0",
								X"01",X"C0",X"07",X"E0",X"03",X"E0",X"0F",X"C0",
								X"07",X"FE",X"7F",X"C0",X"03",X"FF",X"FF",X"80",
								X"01",X"FF",X"FF",X"00",X"00",X"FF",X"FC",X"00",
								X"00",X"1F",X"F0",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- T
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 29
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"0F",X"FF",X"FF",X"E0",X"0F",X"FF",X"FF",X"E0",
								X"0F",X"FF",X"FF",X"E0",X"0F",X"FF",X"FF",X"E0",
								X"00",X"07",X"C0",X"00",X"00",X"07",X"C0",X"00",
								X"00",X"07",X"C0",X"00",X"00",X"07",X"C0",X"00",
								X"00",X"07",X"C0",X"00",X"00",X"07",X"C0",X"00",
								X"00",X"07",X"C0",X"00",X"00",X"07",X"C0",X"00",
								X"00",X"07",X"C0",X"00",X"00",X"07",X"C0",X"00",
								X"00",X"07",X"C0",X"00",X"00",X"07",X"C0",X"00",
								X"00",X"07",X"C0",X"00",X"00",X"07",X"C0",X"00",
								X"00",X"07",X"C0",X"00",X"00",X"07",X"C0",X"00",
								X"00",X"07",X"C0",X"00",X"00",X"07",X"C0",X"00",
								X"00",X"07",X"C0",X"00",X"00",X"07",X"C0",X"00",
								X"00",X"07",X"C0",X"00",X"00",X"07",X"C0",X"00",
								X"00",X"07",X"C0",X"00",X"00",X"07",X"C0",X"00",
								X"00",X"07",X"C0",X"00",X"00",X"07",X"C0",X"00",
								X"00",X"07",X"C0",X"00",X"00",X"07",X"C0",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- U
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 30
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"07",X"E0",X"03",X"E0",X"07",X"C0",X"03",X"E0",
								X"07",X"C0",X"03",X"E0",X"07",X"C0",X"03",X"E0",
								X"07",X"C0",X"03",X"E0",X"07",X"C0",X"03",X"E0",
								X"07",X"C0",X"03",X"E0",X"07",X"C0",X"03",X"E0",
								X"07",X"C0",X"03",X"E0",X"07",X"C0",X"03",X"E0",
								X"07",X"C0",X"03",X"E0",X"07",X"C0",X"03",X"E0",
								X"07",X"C0",X"03",X"E0",X"07",X"C0",X"03",X"E0",
								X"07",X"C0",X"03",X"E0",X"07",X"C0",X"03",X"E0",
								X"07",X"C0",X"03",X"E0",X"07",X"C0",X"03",X"E0",
								X"07",X"C0",X"03",X"E0",X"07",X"C0",X"03",X"E0",
								X"07",X"C0",X"03",X"E0",X"07",X"C0",X"03",X"E0",
								X"07",X"C0",X"03",X"E0",X"07",X"C0",X"03",X"E0",
								X"07",X"E0",X"03",X"E0",X"03",X"E0",X"07",X"C0",
								X"03",X"E0",X"07",X"C0",X"03",X"F0",X"0F",X"C0",
								X"01",X"FC",X"3F",X"80",X"00",X"FF",X"FF",X"00",
								X"00",X"7F",X"FE",X"00",X"00",X"3F",X"FC",X"00",
								X"00",X"0F",X"F0",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- V
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 31
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"0F",X"80",X"01",X"F0",
								X"0F",X"C0",X"01",X"F0",X"07",X"C0",X"01",X"E0",
								X"07",X"C0",X"03",X"E0",X"07",X"E0",X"03",X"E0",
								X"03",X"E0",X"03",X"C0",X"03",X"E0",X"07",X"C0",
								X"03",X"F0",X"07",X"C0",X"01",X"F0",X"07",X"C0",
								X"01",X"F0",X"0F",X"80",X"01",X"F0",X"0F",X"80",
								X"00",X"F8",X"0F",X"80",X"00",X"F8",X"0F",X"00",
								X"00",X"F8",X"1F",X"00",X"00",X"7C",X"1F",X"00",
								X"00",X"7C",X"1E",X"00",X"00",X"7C",X"3E",X"00",
								X"00",X"3E",X"3E",X"00",X"00",X"3E",X"3C",X"00",
								X"00",X"3E",X"7C",X"00",X"00",X"1F",X"7C",X"00",
								X"00",X"1F",X"78",X"00",X"00",X"1F",X"78",X"00",
								X"00",X"0F",X"F8",X"00",X"00",X"0F",X"F0",X"00",
								X"00",X"0F",X"F0",X"00",X"00",X"07",X"F0",X"00",
								X"00",X"07",X"E0",X"00",X"00",X"07",X"E0",X"00",
								X"00",X"03",X"E0",X"00",X"00",X"03",X"C0",X"00",
								X"00",X"03",X"C0",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- W
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 32
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"0F",X"00",X"00",X"F8",X"0F",X"00",X"00",X"F0",
								X"0F",X"01",X"C0",X"F0",X"0F",X"81",X"C0",X"F0",
								X"0F",X"81",X"C0",X"F0",X"0F",X"83",X"E0",X"F0",
								X"07",X"83",X"E0",X"F0",X"07",X"83",X"E0",X"F0",
								X"07",X"83",X"E1",X"E0",X"07",X"87",X"F1",X"E0",
								X"07",X"C7",X"F1",X"E0",X"07",X"C7",X"F1",X"E0",
								X"07",X"C7",X"F1",X"E0",X"03",X"CF",X"79",X"E0",
								X"03",X"CF",X"79",X"E0",X"03",X"CE",X"79",X"C0",
								X"03",X"CE",X"79",X"C0",X"03",X"CE",X"3D",X"C0",
								X"03",X"FE",X"3F",X"C0",X"03",X"FC",X"3F",X"C0",
								X"01",X"FC",X"3F",X"C0",X"01",X"FC",X"1F",X"C0",
								X"01",X"FC",X"1F",X"80",X"01",X"F8",X"1F",X"80",
								X"01",X"F8",X"1F",X"80",X"01",X"F8",X"0F",X"80",
								X"01",X"F8",X"0F",X"80",X"00",X"F0",X"0F",X"80",
								X"00",X"F0",X"0F",X"80",X"00",X"F0",X"07",X"00",
								X"00",X"F0",X"07",X"00",X"00",X"E0",X"07",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- X
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 33
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"07",X"C0",X"03",X"E0",X"03",X"E0",X"07",X"C0",
								X"03",X"E0",X"07",X"C0",X"01",X"F0",X"0F",X"80",
								X"01",X"F8",X"1F",X"80",X"00",X"F8",X"1F",X"00",
								X"00",X"FC",X"3F",X"00",X"00",X"7C",X"3E",X"00",
								X"00",X"7E",X"7E",X"00",X"00",X"3E",X"7C",X"00",
								X"00",X"1F",X"FC",X"00",X"00",X"1F",X"F8",X"00",
								X"00",X"0F",X"F8",X"00",X"00",X"0F",X"F0",X"00",
								X"00",X"07",X"F0",X"00",X"00",X"07",X"E0",X"00",
								X"00",X"07",X"E0",X"00",X"00",X"0F",X"F0",X"00",
								X"00",X"0F",X"F0",X"00",X"00",X"1F",X"F8",X"00",
								X"00",X"1F",X"FC",X"00",X"00",X"3F",X"7C",X"00",
								X"00",X"3E",X"7E",X"00",X"00",X"7E",X"3E",X"00",
								X"00",X"7C",X"3F",X"00",X"00",X"F8",X"1F",X"00",
								X"00",X"F8",X"1F",X"80",X"01",X"F0",X"0F",X"80",
								X"01",X"F0",X"0F",X"C0",X"03",X"E0",X"07",X"E0",
								X"07",X"E0",X"03",X"E0",X"07",X"C0",X"03",X"F0",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- Y
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 34
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"0F",X"C0",X"01",X"F0",X"07",X"C0",X"03",X"E0",
								X"07",X"E0",X"03",X"E0",X"03",X"E0",X"07",X"C0",
								X"03",X"F0",X"07",X"C0",X"01",X"F0",X"0F",X"C0",
								X"01",X"F8",X"0F",X"80",X"00",X"F8",X"0F",X"80",
								X"00",X"FC",X"1F",X"00",X"00",X"7C",X"1F",X"00",
								X"00",X"7E",X"3E",X"00",X"00",X"3E",X"3E",X"00",
								X"00",X"3F",X"7C",X"00",X"00",X"1F",X"7C",X"00",
								X"00",X"1F",X"F8",X"00",X"00",X"0F",X"F8",X"00",
								X"00",X"0F",X"F0",X"00",X"00",X"07",X"F0",X"00",
								X"00",X"07",X"E0",X"00",X"00",X"03",X"E0",X"00",
								X"00",X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",
								X"00",X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",
								X"00",X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",
								X"00",X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",
								X"00",X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",
								X"00",X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- Z
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 35
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"03",X"FF",X"FF",X"E0",X"03",X"FF",X"FF",X"E0",
								X"03",X"FF",X"FF",X"E0",X"03",X"FF",X"FF",X"E0",
								X"00",X"00",X"07",X"C0",X"00",X"00",X"0F",X"80",
								X"00",X"00",X"1F",X"80",X"00",X"00",X"1F",X"00",
								X"00",X"00",X"3F",X"00",X"00",X"00",X"7E",X"00",
								X"00",X"00",X"7C",X"00",X"00",X"00",X"FC",X"00",
								X"00",X"01",X"F8",X"00",X"00",X"01",X"F0",X"00",
								X"00",X"03",X"F0",X"00",X"00",X"03",X"E0",X"00",
								X"00",X"07",X"E0",X"00",X"00",X"0F",X"C0",X"00",
								X"00",X"0F",X"80",X"00",X"00",X"1F",X"80",X"00",
								X"00",X"3F",X"00",X"00",X"00",X"3E",X"00",X"00",
								X"00",X"7E",X"00",X"00",X"00",X"FC",X"00",X"00",
								X"00",X"FC",X"00",X"00",X"01",X"F8",X"00",X"00",
								X"01",X"F0",X"00",X"00",X"03",X"F0",X"00",X"10",
								X"07",X"FF",X"FF",X"F0",X"07",X"FF",X"FF",X"F0",
								X"07",X"FF",X"FF",X"F0",X"07",X"FF",X"FF",X"F0",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- a
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 36
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"0F",X"F0",X"00",
								X"00",X"7F",X"FC",X"00",X"00",X"FF",X"FE",X"00",
								X"03",X"FF",X"FF",X"00",X"01",X"F8",X"3F",X"80",
								X"00",X"E0",X"0F",X"80",X"00",X"00",X"0F",X"C0",
								X"00",X"00",X"07",X"C0",X"00",X"00",X"07",X"C0",
								X"00",X"01",X"FF",X"C0",X"00",X"1F",X"FF",X"C0",
								X"00",X"7F",X"FF",X"C0",X"00",X"FF",X"FF",X"C0",
								X"01",X"FC",X"07",X"C0",X"03",X"F0",X"07",X"C0",
								X"03",X"E0",X"07",X"C0",X"07",X"C0",X"07",X"C0",
								X"07",X"C0",X"0F",X"C0",X"07",X"C0",X"0F",X"C0",
								X"07",X"E0",X"1F",X"C0",X"07",X"F0",X"7F",X"C0",
								X"03",X"FF",X"FF",X"C0",X"01",X"FF",X"F7",X"C0",
								X"00",X"FF",X"E7",X"C0",X"00",X"3F",X"87",X"C0",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- b
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 37
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E1",X"F8",X"00",
								X"03",X"E7",X"FE",X"00",X"03",X"EF",X"FF",X"00",
								X"03",X"FF",X"FF",X"80",X"03",X"FC",X"1F",X"C0",
								X"03",X"F8",X"0F",X"C0",X"03",X"F0",X"07",X"C0",
								X"03",X"F0",X"07",X"E0",X"03",X"E0",X"03",X"E0",
								X"03",X"E0",X"03",X"E0",X"03",X"E0",X"03",X"E0",
								X"03",X"E0",X"03",X"E0",X"03",X"E0",X"03",X"E0",
								X"03",X"E0",X"03",X"E0",X"03",X"E0",X"03",X"E0",
								X"03",X"E0",X"03",X"E0",X"03",X"E0",X"03",X"E0",
								X"03",X"F0",X"07",X"E0",X"03",X"F0",X"07",X"C0",
								X"03",X"F8",X"0F",X"C0",X"03",X"FE",X"3F",X"80",
								X"03",X"FF",X"FF",X"80",X"03",X"DF",X"FF",X"00",
								X"03",X"CF",X"FC",X"00",X"03",X"C3",X"F0",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- c
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 38
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"03",X"F8",X"00",
								X"00",X"0F",X"FF",X"00",X"00",X"3F",X"FF",X"80",
								X"00",X"7F",X"FF",X"C0",X"00",X"FF",X"0F",X"E0",
								X"01",X"FC",X"03",X"C0",X"01",X"F8",X"01",X"80",
								X"03",X"F0",X"01",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"07",X"E0",X"00",X"00",
								X"07",X"E0",X"00",X"00",X"07",X"E0",X"00",X"00",
								X"07",X"E0",X"00",X"00",X"07",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"F0",X"00",X"00",X"01",X"F8",X"01",X"80",
								X"01",X"FC",X"03",X"80",X"00",X"FF",X"1F",X"C0",
								X"00",X"7F",X"FF",X"C0",X"00",X"3F",X"FF",X"80",
								X"00",X"1F",X"FF",X"00",X"00",X"03",X"F8",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- d
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 39
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"E0",
								X"00",X"00",X"07",X"C0",X"00",X"00",X"07",X"C0",
								X"00",X"00",X"07",X"C0",X"00",X"00",X"07",X"C0",
								X"00",X"00",X"07",X"C0",X"00",X"00",X"07",X"C0",
								X"00",X"00",X"07",X"C0",X"00",X"00",X"07",X"C0",
								X"00",X"00",X"07",X"C0",X"00",X"0F",X"C7",X"C0",
								X"00",X"3F",X"F7",X"C0",X"00",X"FF",X"FF",X"C0",
								X"00",X"FF",X"FF",X"C0",X"01",X"F8",X"3F",X"C0",
								X"03",X"F0",X"1F",X"C0",X"03",X"E0",X"0F",X"C0",
								X"07",X"E0",X"0F",X"C0",X"07",X"C0",X"07",X"C0",
								X"07",X"C0",X"07",X"C0",X"07",X"C0",X"07",X"C0",
								X"07",X"C0",X"07",X"C0",X"07",X"C0",X"07",X"C0",
								X"07",X"C0",X"07",X"C0",X"07",X"C0",X"07",X"C0",
								X"07",X"C0",X"07",X"C0",X"07",X"E0",X"07",X"C0",
								X"03",X"E0",X"0F",X"C0",X"03",X"F0",X"0F",X"C0",
								X"03",X"F8",X"1F",X"C0",X"01",X"FC",X"7F",X"C0",
								X"00",X"FF",X"FF",X"C0",X"00",X"7F",X"F7",X"C0",
								X"00",X"3F",X"E7",X"C0",X"00",X"0F",X"C7",X"E0",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- e
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 40
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"07",X"F0",X"00",
								X"00",X"1F",X"FC",X"00",X"00",X"7F",X"FE",X"00",
								X"00",X"FF",X"FF",X"00",X"00",X"FC",X"1F",X"80",
								X"01",X"F0",X"0F",X"80",X"03",X"F0",X"07",X"C0",
								X"03",X"E0",X"07",X"C0",X"03",X"E0",X"07",X"C0",
								X"07",X"C0",X"07",X"C0",X"07",X"FF",X"FF",X"E0",
								X"07",X"FF",X"FF",X"E0",X"07",X"FF",X"FF",X"E0",
								X"07",X"FF",X"FF",X"E0",X"07",X"C0",X"00",X"00",
								X"07",X"C0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"F0",X"00",X"00",
								X"01",X"F8",X"03",X"00",X"01",X"FE",X"0F",X"80",
								X"00",X"FF",X"FF",X"C0",X"00",X"7F",X"FF",X"80",
								X"00",X"1F",X"FE",X"00",X"00",X"07",X"F8",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- f
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 41
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"00",
								X"00",X"01",X"FF",X"C0",X"00",X"07",X"FF",X"E0",
								X"00",X"0F",X"FF",X"F0",X"00",X"0F",X"C1",X"E0",
								X"00",X"1F",X"80",X"E0",X"00",X"1F",X"00",X"40",
								X"00",X"1F",X"00",X"00",X"00",X"1F",X"00",X"00",
								X"00",X"1F",X"00",X"00",X"00",X"1F",X"00",X"00",
								X"07",X"FF",X"FE",X"00",X"07",X"FF",X"FE",X"00",
								X"07",X"FF",X"FE",X"00",X"07",X"FF",X"FE",X"00",
								X"00",X"1F",X"00",X"00",X"00",X"1F",X"00",X"00",
								X"00",X"1F",X"00",X"00",X"00",X"1F",X"00",X"00",
								X"00",X"1F",X"00",X"00",X"00",X"1F",X"00",X"00",
								X"00",X"1F",X"00",X"00",X"00",X"1F",X"00",X"00",
								X"00",X"1F",X"00",X"00",X"00",X"1F",X"00",X"00",
								X"00",X"1F",X"00",X"00",X"00",X"1F",X"00",X"00",
								X"00",X"1F",X"00",X"00",X"00",X"1F",X"00",X"00",
								X"00",X"1F",X"00",X"00",X"00",X"1F",X"00",X"00",
								X"00",X"1F",X"00",X"00",X"00",X"1F",X"00",X"00",
								X"00",X"1F",X"00",X"00",X"00",X"1F",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- g
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 42
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"0F",X"C0",X"F0",X"00",X"3F",X"F7",X"F0",
								X"00",X"7F",X"FF",X"F0",X"00",X"FF",X"FF",X"F0",
								X"01",X"F8",X"7E",X"00",X"01",X"F0",X"3E",X"00",
								X"03",X"E0",X"1E",X"00",X"03",X"E0",X"1F",X"00",
								X"03",X"C0",X"1F",X"00",X"03",X"E0",X"1F",X"00",
								X"03",X"E0",X"1E",X"00",X"01",X"F0",X"3E",X"00",
								X"01",X"F8",X"7E",X"00",X"00",X"FF",X"FC",X"00",
								X"00",X"7F",X"F8",X"00",X"00",X"FF",X"F0",X"00",
								X"01",X"EF",X"C0",X"00",X"01",X"C0",X"00",X"00",
								X"03",X"C0",X"00",X"00",X"03",X"F0",X"00",X"00",
								X"03",X"FF",X"F8",X"00",X"01",X"FF",X"FF",X"00",
								X"00",X"FF",X"FF",X"80",X"01",X"FF",X"FF",X"C0",
								X"03",X"C0",X"3F",X"C0",X"07",X"80",X"03",X"E0",
								X"07",X"80",X"03",X"E0",X"07",X"80",X"03",X"E0",
								X"07",X"80",X"03",X"C0",X"07",X"E0",X"0F",X"C0",
								X"07",X"FF",X"FF",X"80",X"03",X"FF",X"FF",X"00",
								X"00",X"FF",X"FE",X"00",X"00",X"3F",X"F0",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- h
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 43
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"03",X"F0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"F8",X"00",
								X"03",X"E3",X"FE",X"00",X"03",X"E7",X"FF",X"00",
								X"03",X"EF",X"FF",X"80",X"03",X"FE",X"1F",X"80",
								X"03",X"FC",X"0F",X"C0",X"03",X"F8",X"07",X"C0",
								X"03",X"F0",X"07",X"C0",X"03",X"F0",X"07",X"C0",
								X"03",X"E0",X"07",X"C0",X"03",X"E0",X"07",X"C0",
								X"03",X"E0",X"07",X"C0",X"03",X"E0",X"07",X"C0",
								X"03",X"E0",X"07",X"C0",X"03",X"E0",X"07",X"C0",
								X"03",X"E0",X"07",X"C0",X"03",X"E0",X"07",X"C0",
								X"03",X"E0",X"07",X"C0",X"03",X"E0",X"07",X"C0",
								X"03",X"E0",X"07",X"C0",X"03",X"E0",X"07",X"C0",
								X"03",X"E0",X"07",X"C0",X"03",X"E0",X"07",X"C0",
								X"03",X"E0",X"07",X"C0",X"03",X"E0",X"07",X"C0",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- i
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 44
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"07",X"C0",X"00",X"00",X"07",X"E0",X"00",
								X"00",X"07",X"E0",X"00",X"00",X"07",X"E0",X"00",
								X"00",X"07",X"E0",X"00",X"00",X"03",X"C0",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"FF",X"E0",X"00",X"00",X"FF",X"E0",X"00",
								X"00",X"FF",X"E0",X"00",X"00",X"FF",X"E0",X"00",
								X"00",X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",
								X"00",X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",
								X"00",X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",
								X"00",X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",
								X"00",X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",
								X"00",X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",
								X"00",X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",
								X"00",X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",
								X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",
								X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- j
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 45
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"7C",X"00",
								X"00",X"00",X"FE",X"00",X"00",X"00",X"FE",X"00",
								X"00",X"00",X"FE",X"00",X"00",X"00",X"7C",X"00",
								X"00",X"00",X"38",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"7F",X"FE",X"00",X"00",X"7F",X"FE",X"00",
								X"00",X"7F",X"FE",X"00",X"00",X"7F",X"FE",X"00",
								X"00",X"00",X"7E",X"00",X"00",X"00",X"7E",X"00",
								X"00",X"00",X"7E",X"00",X"00",X"00",X"7E",X"00",
								X"00",X"00",X"7E",X"00",X"00",X"00",X"7E",X"00",
								X"00",X"00",X"7E",X"00",X"00",X"00",X"7E",X"00",
								X"00",X"00",X"7E",X"00",X"00",X"00",X"7E",X"00",
								X"00",X"00",X"7E",X"00",X"00",X"00",X"7E",X"00",
								X"00",X"00",X"7E",X"00",X"00",X"00",X"7E",X"00",
								X"00",X"00",X"7E",X"00",X"00",X"00",X"7E",X"00",
								X"00",X"00",X"7E",X"00",X"00",X"00",X"7E",X"00",
								X"00",X"00",X"7E",X"00",X"00",X"00",X"7E",X"00",
								X"00",X"00",X"7E",X"00",X"00",X"80",X"7C",X"00",
								X"01",X"80",X"7C",X"00",X"03",X"C0",X"FC",X"00",
								X"03",X"F3",X"F8",X"00",X"07",X"FF",X"F8",X"00",
								X"03",X"FF",X"F0",X"00",X"01",X"FF",X"C0",X"00",
								X"00",X"3F",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- k
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 46
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"03",X"F0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"0F",X"C0",X"03",X"E0",X"1F",X"80",
								X"03",X"E0",X"3F",X"00",X"03",X"E0",X"7E",X"00",
								X"03",X"E0",X"FC",X"00",X"03",X"E1",X"F8",X"00",
								X"03",X"E3",X"F0",X"00",X"03",X"E7",X"E0",X"00",
								X"03",X"EF",X"C0",X"00",X"03",X"FF",X"80",X"00",
								X"03",X"FF",X"C0",X"00",X"03",X"FF",X"E0",X"00",
								X"03",X"FF",X"F0",X"00",X"03",X"FB",X"F0",X"00",
								X"03",X"F1",X"F8",X"00",X"03",X"E0",X"FC",X"00",
								X"03",X"E0",X"FE",X"00",X"03",X"E0",X"7E",X"00",
								X"03",X"E0",X"3F",X"00",X"03",X"E0",X"1F",X"80",
								X"03",X"E0",X"1F",X"C0",X"03",X"E0",X"0F",X"C0",
								X"03",X"E0",X"07",X"E0",X"03",X"E0",X"03",X"F0",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- l
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 47
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"01",X"FF",X"E0",X"00",
								X"01",X"FF",X"E0",X"00",X"01",X"FF",X"E0",X"00",
								X"01",X"FF",X"E0",X"00",X"00",X"07",X"E0",X"00",
								X"00",X"07",X"E0",X"00",X"00",X"07",X"E0",X"00",
								X"00",X"07",X"E0",X"00",X"00",X"07",X"E0",X"00",
								X"00",X"07",X"E0",X"00",X"00",X"07",X"E0",X"00",
								X"00",X"07",X"E0",X"00",X"00",X"07",X"E0",X"00",
								X"00",X"07",X"E0",X"00",X"00",X"07",X"E0",X"00",
								X"00",X"07",X"E0",X"00",X"00",X"07",X"E0",X"00",
								X"00",X"07",X"E0",X"00",X"00",X"07",X"E0",X"00",
								X"00",X"07",X"E0",X"00",X"00",X"07",X"E0",X"00",
								X"00",X"07",X"E0",X"00",X"00",X"07",X"E0",X"00",
								X"00",X"07",X"E0",X"00",X"00",X"07",X"E0",X"00",
								X"00",X"07",X"E0",X"00",X"00",X"07",X"E0",X"00",
								X"00",X"07",X"E0",X"00",X"00",X"07",X"E0",X"00",
								X"00",X"07",X"E0",X"00",X"00",X"07",X"E0",X"00",
								X"01",X"FF",X"FF",X"80",X"01",X"FF",X"FF",X"80",
								X"01",X"FF",X"FF",X"80",X"01",X"FF",X"FF",X"80",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- m
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 48
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"80",
								X"07",X"BF",X"9F",X"C0",X"07",X"FF",X"BF",X"E0",
								X"07",X"FF",X"FF",X"E0",X"07",X"E7",X"F1",X"F0",
								X"07",X"C3",X"E1",X"F0",X"07",X"C3",X"E1",X"F0",
								X"07",X"83",X"E1",X"F0",X"07",X"83",X"C1",X"F0",
								X"07",X"83",X"C1",X"F0",X"07",X"83",X"C1",X"F0",
								X"07",X"83",X"C1",X"F0",X"07",X"83",X"C1",X"F0",
								X"07",X"83",X"C1",X"F0",X"07",X"83",X"C1",X"F0",
								X"07",X"83",X"C1",X"F0",X"07",X"83",X"C1",X"F0",
								X"07",X"83",X"C1",X"F0",X"07",X"83",X"C1",X"F0",
								X"07",X"83",X"C1",X"F0",X"07",X"83",X"C1",X"F0",
								X"07",X"83",X"C1",X"F0",X"07",X"83",X"C1",X"F0",
								X"07",X"83",X"C1",X"F0",X"07",X"83",X"C1",X"F0",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- n
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 49
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"00",
								X"03",X"E3",X"FE",X"00",X"03",X"E7",X"FF",X"00",
								X"03",X"EF",X"FF",X"80",X"03",X"FE",X"1F",X"80",
								X"03",X"FC",X"0F",X"C0",X"03",X"F8",X"0F",X"C0",
								X"03",X"F0",X"07",X"C0",X"03",X"F0",X"07",X"C0",
								X"03",X"E0",X"07",X"C0",X"03",X"E0",X"07",X"C0",
								X"03",X"E0",X"07",X"C0",X"03",X"E0",X"07",X"C0",
								X"03",X"E0",X"07",X"C0",X"03",X"E0",X"07",X"C0",
								X"03",X"E0",X"07",X"C0",X"03",X"E0",X"07",X"C0",
								X"03",X"E0",X"07",X"C0",X"03",X"E0",X"07",X"C0",
								X"03",X"E0",X"07",X"C0",X"03",X"E0",X"07",X"C0",
								X"03",X"E0",X"07",X"C0",X"03",X"E0",X"07",X"C0",
								X"03",X"E0",X"07",X"C0",X"03",X"E0",X"07",X"C0",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- o
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 50
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"07",X"E0",X"00",
								X"00",X"3F",X"FC",X"00",X"00",X"7F",X"FE",X"00",
								X"00",X"FF",X"FF",X"00",X"01",X"FC",X"3F",X"80",
								X"03",X"F0",X"0F",X"C0",X"03",X"F0",X"0F",X"C0",
								X"07",X"E0",X"07",X"E0",X"07",X"E0",X"07",X"E0",
								X"07",X"C0",X"03",X"E0",X"07",X"C0",X"03",X"E0",
								X"07",X"C0",X"03",X"E0",X"07",X"C0",X"03",X"E0",
								X"07",X"C0",X"03",X"E0",X"07",X"C0",X"03",X"E0",
								X"07",X"C0",X"03",X"E0",X"07",X"E0",X"07",X"E0",
								X"07",X"E0",X"07",X"E0",X"03",X"F0",X"0F",X"C0",
								X"03",X"F8",X"1F",X"C0",X"01",X"FC",X"3F",X"80",
								X"00",X"FF",X"FF",X"00",X"00",X"7F",X"FE",X"00",
								X"00",X"3F",X"FC",X"00",X"00",X"0F",X"E0",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- p
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 51
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"01",X"F8",X"00",
								X"03",X"E7",X"FE",X"00",X"03",X"EF",X"FF",X"00",
								X"03",X"FF",X"FF",X"80",X"03",X"FE",X"3F",X"C0",
								X"03",X"F8",X"0F",X"C0",X"03",X"F0",X"07",X"E0",
								X"03",X"F0",X"07",X"E0",X"03",X"E0",X"03",X"E0",
								X"03",X"E0",X"03",X"E0",X"03",X"E0",X"03",X"E0",
								X"03",X"E0",X"03",X"E0",X"03",X"E0",X"03",X"E0",
								X"03",X"E0",X"03",X"E0",X"03",X"E0",X"03",X"E0",
								X"03",X"E0",X"03",X"E0",X"03",X"E0",X"03",X"E0",
								X"03",X"F0",X"07",X"E0",X"03",X"F0",X"07",X"C0",
								X"03",X"F8",X"0F",X"C0",X"03",X"FC",X"3F",X"80",
								X"03",X"FF",X"FF",X"80",X"03",X"FF",X"FF",X"00",
								X"03",X"E7",X"FE",X"00",X"03",X"E3",X"F8",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"E0",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- q
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 52
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"0F",X"C0",X"00",
								X"00",X"3F",X"F7",X"C0",X"00",X"FF",X"FF",X"C0",
								X"01",X"FF",X"FF",X"C0",X"01",X"FC",X"3F",X"C0",
								X"03",X"F0",X"1F",X"C0",X"03",X"E0",X"0F",X"C0",
								X"07",X"E0",X"07",X"C0",X"07",X"C0",X"07",X"C0",
								X"07",X"C0",X"07",X"C0",X"07",X"C0",X"07",X"C0",
								X"07",X"C0",X"07",X"C0",X"07",X"C0",X"07",X"C0",
								X"07",X"C0",X"07",X"C0",X"07",X"C0",X"07",X"C0",
								X"07",X"C0",X"07",X"C0",X"07",X"C0",X"07",X"C0",
								X"07",X"E0",X"0F",X"C0",X"03",X"E0",X"0F",X"C0",
								X"03",X"F0",X"1F",X"C0",X"01",X"FC",X"7F",X"C0",
								X"01",X"FF",X"FF",X"C0",X"00",X"FF",X"FF",X"C0",
								X"00",X"3F",X"F7",X"C0",X"00",X"0F",X"C7",X"C0",
								X"00",X"00",X"07",X"C0",X"00",X"00",X"07",X"C0",
								X"00",X"00",X"07",X"C0",X"00",X"00",X"07",X"C0",
								X"00",X"00",X"07",X"C0",X"00",X"00",X"07",X"C0",
								X"00",X"00",X"07",X"C0",X"00",X"00",X"07",X"C0",
								X"00",X"00",X"07",X"C0"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- r
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 53
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"00",
								X"00",X"FC",X"FF",X"C0",X"00",X"FD",X"FF",X"E0",
								X"00",X"FB",X"FF",X"E0",X"00",X"FF",X"E7",X"C0",
								X"00",X"FF",X"01",X"C0",X"00",X"FE",X"00",X"80",
								X"00",X"FC",X"00",X"00",X"00",X"FC",X"00",X"00",
								X"00",X"FC",X"00",X"00",X"00",X"FC",X"00",X"00",
								X"00",X"F8",X"00",X"00",X"00",X"F8",X"00",X"00",
								X"00",X"F8",X"00",X"00",X"00",X"F8",X"00",X"00",
								X"00",X"F8",X"00",X"00",X"00",X"F8",X"00",X"00",
								X"00",X"F8",X"00",X"00",X"00",X"F8",X"00",X"00",
								X"00",X"F8",X"00",X"00",X"00",X"F8",X"00",X"00",
								X"00",X"F8",X"00",X"00",X"00",X"F8",X"00",X"00",
								X"00",X"F8",X"00",X"00",X"00",X"F8",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- s
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 54
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"0F",X"F0",X"00",
								X"00",X"3F",X"FE",X"00",X"00",X"7F",X"FF",X"00",
								X"00",X"FF",X"FF",X"C0",X"01",X"F8",X"1F",X"80",
								X"01",X"F0",X"07",X"80",X"01",X"F0",X"03",X"00",
								X"01",X"F0",X"00",X"00",X"01",X"F8",X"00",X"00",
								X"00",X"FF",X"00",X"00",X"00",X"7F",X"E0",X"00",
								X"00",X"3F",X"FC",X"00",X"00",X"0F",X"FF",X"00",
								X"00",X"03",X"FF",X"80",X"00",X"00",X"7F",X"C0",
								X"00",X"00",X"0F",X"C0",X"00",X"80",X"07",X"C0",
								X"00",X"80",X"07",X"C0",X"01",X"C0",X"07",X"C0",
								X"03",X"E0",X"07",X"C0",X"03",X"F8",X"1F",X"C0",
								X"03",X"FF",X"FF",X"80",X"01",X"FF",X"FF",X"00",
								X"00",X"7F",X"FE",X"00",X"00",X"0F",X"F0",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- t
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 55
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"07",X"80",X"00",
								X"00",X"0F",X"80",X"00",X"00",X"1F",X"80",X"00",
								X"00",X"1F",X"80",X"00",X"00",X"1F",X"80",X"00",
								X"00",X"1F",X"80",X"00",X"00",X"1F",X"00",X"00",
								X"03",X"FF",X"FF",X"00",X"03",X"FF",X"FF",X"00",
								X"03",X"FF",X"FF",X"00",X"03",X"FF",X"FF",X"00",
								X"00",X"1F",X"00",X"00",X"00",X"1F",X"00",X"00",
								X"00",X"1F",X"00",X"00",X"00",X"1F",X"00",X"00",
								X"00",X"1F",X"00",X"00",X"00",X"1F",X"00",X"00",
								X"00",X"1F",X"00",X"00",X"00",X"1F",X"00",X"00",
								X"00",X"1F",X"00",X"00",X"00",X"1F",X"00",X"00",
								X"00",X"1F",X"00",X"00",X"00",X"1F",X"00",X"00",
								X"00",X"1F",X"00",X"00",X"00",X"1F",X"80",X"00",
								X"00",X"1F",X"80",X"C0",X"00",X"0F",X"C3",X"C0",
								X"00",X"0F",X"FF",X"C0",X"00",X"07",X"FF",X"C0",
								X"00",X"03",X"FF",X"80",X"00",X"01",X"FC",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- u
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 56
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"03",X"E0",X"07",X"C0",X"03",X"E0",X"07",X"C0",
								X"03",X"E0",X"07",X"C0",X"03",X"E0",X"07",X"C0",
								X"03",X"E0",X"07",X"C0",X"03",X"E0",X"07",X"C0",
								X"03",X"E0",X"07",X"C0",X"03",X"E0",X"07",X"C0",
								X"03",X"E0",X"07",X"C0",X"03",X"E0",X"07",X"C0",
								X"03",X"E0",X"07",X"C0",X"03",X"E0",X"07",X"C0",
								X"03",X"E0",X"07",X"C0",X"03",X"E0",X"07",X"C0",
								X"03",X"E0",X"07",X"C0",X"03",X"E0",X"0F",X"C0",
								X"03",X"E0",X"0F",X"C0",X"03",X"F0",X"0F",X"C0",
								X"03",X"F0",X"1F",X"C0",X"01",X"FC",X"7F",X"C0",
								X"01",X"FF",X"FF",X"C0",X"00",X"FF",X"F7",X"C0",
								X"00",X"7F",X"E7",X"C0",X"00",X"1F",X"87",X"C0",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- v
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 57
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"07",X"C0",X"03",X"E0",X"07",X"E0",X"03",X"E0",
								X"03",X"E0",X"03",X"C0",X"03",X"E0",X"03",X"C0",
								X"03",X"F0",X"07",X"C0",X"01",X"F0",X"07",X"C0",
								X"01",X"F0",X"07",X"80",X"00",X"F8",X"0F",X"80",
								X"00",X"F8",X"0F",X"00",X"00",X"FC",X"0F",X"00",
								X"00",X"7C",X"1F",X"00",X"00",X"7C",X"1E",X"00",
								X"00",X"7E",X"3E",X"00",X"00",X"3E",X"3C",X"00",
								X"00",X"3E",X"7C",X"00",X"00",X"1F",X"7C",X"00",
								X"00",X"1F",X"78",X"00",X"00",X"1F",X"F8",X"00",
								X"00",X"0F",X"F0",X"00",X"00",X"0F",X"F0",X"00",
								X"00",X"07",X"E0",X"00",X"00",X"07",X"E0",X"00",
								X"00",X"07",X"E0",X"00",X"00",X"03",X"C0",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- w
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 58
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"0F",X"00",X"00",X"F0",X"0F",X"00",X"00",X"F0",
								X"0F",X"00",X"00",X"F0",X"0F",X"81",X"C0",X"F0",
								X"0F",X"83",X"C0",X"F0",X"07",X"83",X"C0",X"F0",
								X"07",X"83",X"E1",X"E0",X"07",X"83",X"E1",X"E0",
								X"07",X"C7",X"E1",X"E0",X"07",X"C7",X"F1",X"E0",
								X"03",X"C7",X"F1",X"E0",X"03",X"C7",X"71",X"E0",
								X"03",X"CF",X"79",X"E0",X"03",X"CE",X"79",X"C0",
								X"03",X"EE",X"7B",X"C0",X"01",X"EE",X"3F",X"C0",
								X"01",X"FE",X"3F",X"C0",X"01",X"FC",X"3F",X"C0",
								X"01",X"FC",X"3F",X"C0",X"01",X"FC",X"1F",X"80",
								X"01",X"FC",X"1F",X"80",X"00",X"F8",X"1F",X"80",
								X"00",X"F8",X"1F",X"80",X"00",X"F8",X"0F",X"80",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- x
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 59
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"07",X"E0",X"07",X"C0",X"03",X"E0",X"0F",X"80",
								X"01",X"F0",X"1F",X"80",X"01",X"F8",X"1F",X"00",
								X"00",X"FC",X"3E",X"00",X"00",X"7C",X"3E",X"00",
								X"00",X"7E",X"7C",X"00",X"00",X"3F",X"F8",X"00",
								X"00",X"1F",X"F8",X"00",X"00",X"1F",X"F0",X"00",
								X"00",X"0F",X"F0",X"00",X"00",X"07",X"E0",X"00",
								X"00",X"07",X"E0",X"00",X"00",X"0F",X"F0",X"00",
								X"00",X"1F",X"F8",X"00",X"00",X"1F",X"F8",X"00",
								X"00",X"3E",X"FC",X"00",X"00",X"7E",X"7E",X"00",
								X"00",X"7C",X"3E",X"00",X"00",X"F8",X"1F",X"00",
								X"01",X"F8",X"1F",X"80",X"03",X"F0",X"0F",X"C0",
								X"03",X"E0",X"07",X"C0",X"07",X"E0",X"07",X"E0",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- y
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 60
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"07",X"C0",X"07",X"C0",X"07",X"E0",X"07",X"C0",
								X"03",X"E0",X"07",X"C0",X"03",X"E0",X"07",X"C0",
								X"01",X"F0",X"07",X"C0",X"01",X"F0",X"0F",X"80",
								X"01",X"F8",X"0F",X"80",X"00",X"F8",X"0F",X"80",
								X"00",X"F8",X"0F",X"00",X"00",X"7C",X"1F",X"00",
								X"00",X"7C",X"1E",X"00",X"00",X"3E",X"1E",X"00",
								X"00",X"3E",X"3E",X"00",X"00",X"3E",X"3C",X"00",
								X"00",X"1F",X"7C",X"00",X"00",X"1F",X"7C",X"00",
								X"00",X"0F",X"F8",X"00",X"00",X"0F",X"F8",X"00",
								X"00",X"0F",X"F0",X"00",X"00",X"07",X"F0",X"00",
								X"00",X"07",X"F0",X"00",X"00",X"03",X"E0",X"00",
								X"00",X"03",X"E0",X"00",X"00",X"03",X"E0",X"00",
								X"00",X"03",X"C0",X"00",X"00",X"03",X"C0",X"00",
								X"00",X"07",X"C0",X"00",X"02",X"0F",X"80",X"00",
								X"07",X"1F",X"80",X"00",X"07",X"FF",X"00",X"00",
								X"0F",X"FE",X"00",X"00",X"07",X"FC",X"00",X"00",
								X"01",X"F0",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- z
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 61
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"03",X"FF",X"FF",X"C0",X"03",X"FF",X"FF",X"C0",
								X"03",X"FF",X"FF",X"C0",X"03",X"FF",X"FF",X"80",
								X"00",X"00",X"1F",X"80",X"00",X"00",X"3F",X"00",
								X"00",X"00",X"7E",X"00",X"00",X"00",X"FC",X"00",
								X"00",X"00",X"F8",X"00",X"00",X"01",X"F0",X"00",
								X"00",X"03",X"F0",X"00",X"00",X"07",X"E0",X"00",
								X"00",X"0F",X"C0",X"00",X"00",X"1F",X"80",X"00",
								X"00",X"1F",X"00",X"00",X"00",X"3E",X"00",X"00",
								X"00",X"7E",X"00",X"00",X"00",X"FC",X"00",X"00",
								X"01",X"F8",X"00",X"00",X"03",X"F0",X"00",X"20",
								X"03",X"FF",X"FF",X"E0",X"07",X"FF",X"FF",X"E0",
								X"07",X"FF",X"FF",X"E0",X"07",X"FF",X"FF",X"E0",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --!
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  --62
								X"00",X"00",X"00",X"00",X"00",X"03",X"C0",X"00",
								X"00",X"03",X"C0",X"00",X"00",X"03",X"C0",X"00",
								X"00",X"03",X"C0",X"00",X"00",X"03",X"C0",X"00",
								X"00",X"03",X"C0",X"00",X"00",X"03",X"C0",X"00",
								X"00",X"03",X"C0",X"00",X"00",X"03",X"C0",X"00",
								X"00",X"03",X"C0",X"00",X"00",X"03",X"C0",X"00",
								X"00",X"03",X"C0",X"00",X"00",X"03",X"C0",X"00",
								X"00",X"03",X"C0",X"00",X"00",X"03",X"80",X"00",
								X"00",X"03",X"80",X"00",X"00",X"03",X"80",X"00",
								X"00",X"03",X"80",X"00",X"00",X"03",X"80",X"00",
								X"00",X"03",X"80",X"00",X"00",X"03",X"80",X"00",
								X"00",X"03",X"80",X"00",X"00",X"03",X"80",X"00",
								X"00",X"03",X"80",X"00",X"00",X"03",X"80",X"00",
								X"00",X"03",X"80",X"00",X"00",X"03",X"80",X"00",
								X"00",X"03",X"80",X"00",X"00",X"03",X"80",X"00",
								X"00",X"03",X"80",X"00",X"00",X"03",X"80",X"00",
								X"00",X"03",X"80",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"01",X"80",X"00",
								X"00",X"07",X"C0",X"00",X"00",X"07",X"C0",X"00",
								X"00",X"07",X"C0",X"00",X"00",X"07",X"C0",X"00",
								X"00",X"07",X"C0",X"00",X"00",X"03",X"80",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --"
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --63
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"78",X"1C",X"00",
								X"00",X"78",X"3E",X"00",X"00",X"78",X"3E",X"00",
								X"00",X"78",X"3E",X"00",X"00",X"78",X"3E",X"00",
								X"00",X"78",X"3E",X"00",X"00",X"78",X"3E",X"00",
								X"00",X"78",X"3E",X"00",X"00",X"78",X"3E",X"00",
								X"00",X"78",X"3E",X"00",X"00",X"78",X"3E",X"00",
								X"00",X"78",X"3E",X"00",X"00",X"78",X"3E",X"00",
								X"00",X"78",X"3E",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --#
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  --64
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"07",X"07",X"00",X"00",X"07",X"07",X"00",
								X"00",X"07",X"06",X"00",X"00",X"06",X"0E",X"00",
								X"00",X"0E",X"0E",X"00",X"00",X"0E",X"0E",X"00",
								X"00",X"0E",X"0E",X"00",X"00",X"0E",X"0C",X"00",
								X"00",X"0C",X"1C",X"00",X"07",X"FF",X"FF",X"F0",
								X"07",X"FF",X"FF",X"F0",X"00",X"3C",X"3C",X"00",
								X"00",X"1C",X"18",X"00",X"00",X"18",X"38",X"00",
								X"00",X"38",X"38",X"00",X"00",X"38",X"38",X"00",
								X"00",X"38",X"38",X"00",X"00",X"30",X"70",X"00",
								X"00",X"78",X"70",X"00",X"1F",X"FF",X"FF",X"C0",
								X"1F",X"FF",X"FF",X"C0",X"00",X"60",X"60",X"00",
								X"00",X"60",X"E0",X"00",X"00",X"E0",X"E0",X"00",
								X"00",X"E0",X"E0",X"00",X"00",X"E0",X"C0",X"00",
								X"00",X"C0",X"C0",X"00",X"01",X"C0",X"C0",X"00",
								X"01",X"C0",X"C0",X"00",X"01",X"C0",X"C0",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --%
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  --65
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"03",X"F0",X"07",X"00",X"07",X"F8",X"06",X"00",
								X"0E",X"1C",X"0C",X"00",X"0C",X"0C",X"1C",X"00",
								X"1C",X"0C",X"18",X"00",X"18",X"0C",X"30",X"00",
								X"18",X"0C",X"70",X"00",X"1C",X"0C",X"60",X"00",
								X"0C",X"0C",X"E0",X"00",X"0C",X"1C",X"C0",X"00",
								X"0E",X"38",X"80",X"00",X"01",X"C1",X"0F",X"80",
								X"00",X"03",X"1F",X"C0",X"00",X"07",X"30",X"60",
								X"00",X"06",X"70",X"70",X"00",X"0E",X"60",X"30",
								X"00",X"0C",X"60",X"30",X"00",X"18",X"60",X"30",
								X"00",X"38",X"60",X"30",X"00",X"30",X"60",X"70",
								X"00",X"60",X"70",X"60",X"00",X"E0",X"38",X"E0",
								X"00",X"C0",X"1F",X"C0",X"00",X"80",X"0F",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --&
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  --66
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"3F",X"00",X"00",
								X"00",X"7F",X"80",X"00",X"00",X"E1",X"C0",X"00",
								X"01",X"C0",X"C0",X"00",X"01",X"C0",X"C0",X"00",
								X"01",X"80",X"C0",X"00",X"01",X"C0",X"C1",X"C0",
								X"00",X"C0",X"C1",X"C0",X"00",X"E1",X"81",X"C0",
								X"00",X"7F",X"01",X"C0",X"00",X"7E",X"01",X"80",
								X"00",X"FF",X"01",X"80",X"03",X"80",X"C3",X"80",
								X"07",X"00",X"E3",X"00",X"06",X"00",X"77",X"00",
								X"0E",X"00",X"7E",X"00",X"0E",X"00",X"3E",X"00",
								X"0E",X"00",X"1C",X"00",X"0E",X"00",X"3C",X"00",
								X"07",X"00",X"7E",X"00",X"07",X"80",X"F7",X"00",
								X"03",X"FF",X"C3",X"F0",X"01",X"FF",X"81",X"F0",
								X"00",X"3E",X"00",X"E0",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --'
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  --67
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",
								X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"00",
								X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"00",
								X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"00",
								X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --(
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  --68
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",
								X"00",X"00",X"80",X"00",X"00",X"01",X"80",X"00",
								X"00",X"01",X"00",X"00",X"00",X"03",X"00",X"00",
								X"00",X"03",X"00",X"00",X"00",X"06",X"00",X"00",
								X"00",X"06",X"00",X"00",X"00",X"0E",X"00",X"00",
								X"00",X"0C",X"00",X"00",X"00",X"0C",X"00",X"00",
								X"00",X"0C",X"00",X"00",X"00",X"0C",X"00",X"00",
								X"00",X"0C",X"00",X"00",X"00",X"0C",X"00",X"00",
								X"00",X"0C",X"00",X"00",X"00",X"0C",X"00",X"00",
								X"00",X"0C",X"00",X"00",X"00",X"0C",X"00",X"00",
								X"00",X"0C",X"00",X"00",X"00",X"0C",X"00",X"00",
								X"00",X"0E",X"00",X"00",X"00",X"06",X"00",X"00",
								X"00",X"06",X"00",X"00",X"00",X"07",X"00",X"00",
								X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"00",
								X"00",X"01",X"00",X"00",X"00",X"01",X"80",X"00",
								X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --)
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  --69
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",
								X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"00",
								X"00",X"01",X"00",X"00",X"00",X"01",X"80",X"00",
								X"00",X"00",X"80",X"00",X"00",X"00",X"C0",X"00",
								X"00",X"00",X"C0",X"00",X"00",X"00",X"C0",X"00",
								X"00",X"00",X"C0",X"00",X"00",X"00",X"E0",X"00",
								X"00",X"00",X"60",X"00",X"00",X"00",X"60",X"00",
								X"00",X"00",X"60",X"00",X"00",X"00",X"60",X"00",
								X"00",X"00",X"60",X"00",X"00",X"00",X"60",X"00",
								X"00",X"00",X"60",X"00",X"00",X"00",X"60",X"00",
								X"00",X"00",X"E0",X"00",X"00",X"00",X"C0",X"00",
								X"00",X"00",X"C0",X"00",X"00",X"00",X"C0",X"00",
								X"00",X"00",X"C0",X"00",X"00",X"00",X"80",X"00",
								X"00",X"01",X"80",X"00",X"00",X"01",X"00",X"00",
								X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"00",
								X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --*
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  --70
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",
								X"00",X"1D",X"38",X"00",X"00",X"0F",X"F0",X"00",
								X"00",X"01",X"80",X"00",X"00",X"03",X"C0",X"00",
								X"00",X"06",X"E0",X"00",X"00",X"0E",X"60",X"00",
								X"00",X"04",X"20",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --+
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  --71
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
								X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",
								X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",
								X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",
								X"00",X"FF",X"FE",X"00",X"00",X"01",X"80",X"00",
								X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",
								X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",
								X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --,
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  --72
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
								X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",
								X"00",X"01",X"00",X"00",X"00",X"03",X"00",X"00",
								X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- -
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  --73
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"0F",X"F0",X"00",
								X"00",X"0F",X"F0",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --.
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  --74
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",
								X"00",X"07",X"00",X"00",X"00",X"07",X"80",X"00",
								X"00",X"07",X"00",X"00",X"00",X"03",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --/
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  --75
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",
								X"00",X"00",X"07",X"80",X"00",X"00",X"07",X"00",
								X"00",X"00",X"0F",X"00",X"00",X"00",X"0E",X"00",
								X"00",X"00",X"1E",X"00",X"00",X"00",X"1E",X"00",
								X"00",X"00",X"1C",X"00",X"00",X"00",X"3C",X"00",
								X"00",X"00",X"38",X"00",X"00",X"00",X"78",X"00",
								X"00",X"00",X"78",X"00",X"00",X"00",X"70",X"00",
								X"00",X"00",X"F0",X"00",X"00",X"00",X"E0",X"00",
								X"00",X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",
								X"00",X"00",X"C0",X"00",X"00",X"01",X"C0",X"00",
								X"00",X"01",X"80",X"00",X"00",X"03",X"80",X"00",
								X"00",X"03",X"00",X"00",X"00",X"07",X"00",X"00",
								X"00",X"07",X"00",X"00",X"00",X"0F",X"00",X"00",
								X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",
								X"00",X"1E",X"00",X"00",X"00",X"1C",X"00",X"00",
								X"00",X"3C",X"00",X"00",X"00",X"38",X"00",X"00",
								X"00",X"38",X"00",X"00",X"00",X"78",X"00",X"00",
								X"00",X"70",X"00",X"00",X"00",X"F0",X"00",X"00",
								X"00",X"E0",X"00",X"00",X"00",X"E0",X"00",X"00",
								X"01",X"E0",X"00",X"00",X"01",X"C0",X"00",X"00",
								X"01",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --:
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  --76
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"03",X"00",X"00",X"00",X"03",X"80",X"00",
								X"00",X"03",X"80",X"00",X"00",X"03",X"00",X"00",
								X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",
								X"00",X"03",X"00",X"00",X"00",X"03",X"80",X"00",
								X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --;
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  --77
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"01",X"00",X"00",X"00",X"03",X"80",X"00",
								X"00",X"03",X"C0",X"00",X"00",X"03",X"C0",X"00",
								X"00",X"01",X"80",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"01",X"80",X"00",
								X"00",X"01",X"80",X"00",X"00",X"03",X"80",X"00",
								X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"00",
								X"00",X"03",X"00",X"00",X"00",X"07",X"00",X"00",
								X"00",X"07",X"00",X"00",X"00",X"07",X"00",X"00",
								X"00",X"06",X"00",X"00",X"00",X"0E",X"00",X"00",
								X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --<
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  --78
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",
								X"00",X"00",X"1F",X"00",X"00",X"00",X"7E",X"00",
								X"00",X"00",X"FC",X"00",X"00",X"01",X"F0",X"00",
								X"00",X"07",X"C0",X"00",X"00",X"1F",X"00",X"00",
								X"00",X"7E",X"00",X"00",X"00",X"FC",X"00",X"00",
								X"03",X"F0",X"00",X"00",X"07",X"E0",X"00",X"00",
								X"01",X"F8",X"00",X"00",X"00",X"7E",X"00",X"00",
								X"00",X"1F",X"00",X"00",X"00",X"07",X"C0",X"00",
								X"00",X"01",X"F0",X"00",X"00",X"00",X"FC",X"00",
								X"00",X"00",X"3E",X"00",X"00",X"00",X"1F",X"00",
								X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --=
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  --79
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"07",X"FF",X"FF",X"C0",X"07",X"FF",X"FF",X"C0",
								X"07",X"FF",X"FF",X"C0",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"07",X"FF",X"FF",X"C0",
								X"07",X"FF",X"FF",X"C0",X"07",X"FF",X"FF",X"C0",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -->
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  --80
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"02",X"00",X"00",X"00",X"03",X"80",X"00",X"00",
								X"03",X"E0",X"00",X"00",X"01",X"F0",X"00",X"00",
								X"00",X"FC",X"00",X"00",X"00",X"3F",X"00",X"00",
								X"00",X"0F",X"80",X"00",X"00",X"03",X"E0",X"00",
								X"00",X"00",X"F0",X"00",X"00",X"00",X"FC",X"00",
								X"00",X"00",X"3F",X"00",X"00",X"00",X"0F",X"80",
								X"00",X"00",X"3F",X"00",X"00",X"00",X"FC",X"00",
								X"00",X"01",X"F0",X"00",X"00",X"0F",X"C0",X"00",
								X"00",X"3F",X"00",X"00",X"00",X"FE",X"00",X"00",
								X"01",X"F8",X"00",X"00",X"03",X"E0",X"00",X"00",
								X"03",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --?
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  --81
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"07",X"E0",X"00",
								X"00",X"3F",X"FC",X"00",X"00",X"7F",X"FE",X"00",
								X"00",X"78",X"3E",X"00",X"00",X"60",X"1F",X"00",
								X"00",X"40",X"0F",X"00",X"00",X"00",X"0F",X"00",
								X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",
								X"00",X"00",X"0F",X"00",X"00",X"00",X"1E",X"00",
								X"00",X"00",X"1E",X"00",X"00",X"00",X"3C",X"00",
								X"00",X"00",X"78",X"00",X"00",X"00",X"F0",X"00",
								X"00",X"00",X"E0",X"00",X"00",X"03",X"80",X"00",
								X"00",X"03",X"00",X"00",X"00",X"07",X"00",X"00",
								X"00",X"07",X"00",X"00",X"00",X"07",X"00",X"00",
								X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"03",X"80",X"00",
								X"00",X"03",X"80",X"00",X"00",X"03",X"80",X"00",
								X"00",X"03",X"80",X"00",X"00",X"01",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --deg c
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  --82
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"1F",X"F8",X"00",X"00",X"1F",X"F8",X"00",X"00",
								X"1F",X"F8",X"00",X"00",X"1C",X"38",X"00",X"00",
								X"1C",X"38",X"00",X"00",X"1C",X"38",X"00",X"00",
								X"1C",X"38",X"00",X"00",X"1F",X"F8",X"00",X"00",
								X"1F",X"F8",X"00",X"00",X"1F",X"F8",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"03",X"FF",X"F8",
								X"00",X"07",X"FF",X"F8",X"00",X"07",X"FF",X"F8",
								X"00",X"07",X"00",X"00",X"00",X"07",X"00",X"00",
								X"00",X"07",X"00",X"00",X"00",X"07",X"00",X"00",
								X"00",X"07",X"00",X"00",X"00",X"07",X"00",X"00",
								X"00",X"07",X"00",X"00",X"00",X"07",X"00",X"00",
								X"00",X"07",X"00",X"00",X"00",X"07",X"00",X"00",
								X"00",X"07",X"00",X"00",X"00",X"07",X"00",X"00",
								X"00",X"07",X"FF",X"FC",X"00",X"07",X"FF",X"FC",
								X"00",X"03",X"FF",X"FC",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00")
								);
    --------------------------------------------------------------------------------
	-- 0~9 A~Z a~z
    type rom26x16 is array (0 to 84, 0 to 51) of std_logic_vector(7 downto 0); 
	constant Font26 : rom26x16 :=( -- 26 x 16 / 8 = 52 Bytes (rows x cols = H x W)
								(X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"C0", -- 0
								X"0F",X"E0",X"1E",X"F0",X"3C",X"78",X"38",X"38",  -- 0
								X"38",X"38",X"30",X"78",X"70",X"DC",X"71",X"DC",
								X"73",X"9C",X"73",X"1C",X"76",X"1C",X"3C",X"18",
								X"38",X"38",X"38",X"38",X"38",X"38",X"1E",X"F0",
								X"0F",X"E0",X"07",X"C0",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"80", -- 1
								X"0F",X"80",X"1F",X"80",X"1F",X"80",X"03",X"80",  -- 1
								X"03",X"80",X"03",X"80",X"03",X"80",X"03",X"80",
								X"03",X"80",X"03",X"80",X"03",X"80",X"03",X"80",
								X"03",X"80",X"03",X"80",X"03",X"80",X"03",X"80",
								X"03",X"80",X"03",X"80",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"C0", -- 2
								X"1F",X"F0",X"3F",X"F8",X"78",X"38",X"10",X"38",  -- 2
								X"00",X"38",X"00",X"38",X"00",X"38",X"00",X"78",
								X"00",X"70",X"00",X"E0",X"01",X"E0",X"03",X"C0",
								X"07",X"80",X"0F",X"00",X"1E",X"00",X"3C",X"08",
								X"3F",X"F8",X"3F",X"F8",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"C0", -- 3
								X"1F",X"E0",X"3F",X"F0",X"10",X"70",X"00",X"38",  -- 3
								X"00",X"30",X"00",X"70",X"01",X"E0",X"07",X"C0",
								X"07",X"E0",X"00",X"70",X"00",X"38",X"00",X"38",
								X"00",X"38",X"10",X"38",X"10",X"78",X"3D",X"F0",
								X"3F",X"E0",X"0F",X"C0",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70", -- 4
								X"00",X"F0",X"00",X"F0",X"01",X"F0",X"03",X"F0",  -- 4
								X"03",X"70",X"07",X"70",X"0E",X"70",X"0C",X"70",
								X"1C",X"70",X"38",X"70",X"30",X"70",X"7F",X"FC",
								X"7F",X"FC",X"00",X"70",X"00",X"70",X"00",X"70",
								X"00",X"70",X"00",X"70",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"F8", -- 5
								X"1F",X"F8",X"1C",X"00",X"18",X"00",X"18",X"00",  -- 5
								X"18",X"00",X"1B",X"C0",X"1F",X"F0",X"3E",X"F8",
								X"18",X"38",X"00",X"38",X"00",X"1C",X"00",X"1C",
								X"00",X"1C",X"00",X"38",X"38",X"38",X"3E",X"F8",
								X"1F",X"F0",X"07",X"C0",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"E0", -- 6
								X"07",X"F8",X"0F",X"F0",X"1C",X"10",X"1C",X"00",  -- 6
								X"38",X"00",X"38",X"00",X"3B",X"E0",X"3F",X"F0",
								X"3E",X"78",X"38",X"38",X"38",X"18",X"38",X"18",
								X"38",X"18",X"38",X"38",X"1C",X"38",X"1F",X"F0",
								X"0F",X"F0",X"07",X"C0",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"F8", -- 7
								X"3F",X"F8",X"3F",X"F8",X"00",X"70",X"00",X"70",  -- 7
								X"00",X"70",X"00",X"E0",X"00",X"E0",X"00",X"E0",
								X"01",X"C0",X"01",X"C0",X"03",X"80",X"03",X"80",
								X"03",X"80",X"07",X"80",X"07",X"00",X"07",X"00",
								X"0F",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"C0", -- 8
								X"0F",X"F0",X"1E",X"F0",X"38",X"38",X"38",X"38",  -- 8
								X"38",X"38",X"1C",X"38",X"1E",X"70",X"0F",X"E0",
								X"0F",X"E0",X"1C",X"F0",X"38",X"38",X"38",X"38",
								X"70",X"1C",X"78",X"1C",X"38",X"38",X"3F",X"F8",
								X"1F",X"F0",X"07",X"C0",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"C0", -- 9
								X"0F",X"E0",X"1E",X"F0",X"38",X"38",X"38",X"38",  -- 9
								X"30",X"38",X"30",X"38",X"38",X"18",X"38",X"38",
								X"3E",X"F8",X"1F",X"F8",X"07",X"F8",X"00",X"38",
								X"00",X"38",X"00",X"30",X"10",X"70",X"3D",X"E0",
								X"3F",X"E0",X"0F",X"80",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00", -- A
								X"03",X"80",X"03",X"80",X"03",X"80",X"07",X"C0",  -- 10
								X"07",X"C0",X"06",X"C0",X"0E",X"E0",X"0E",X"E0",
								X"0C",X"60",X"1C",X"70",X"1C",X"70",X"1F",X"F0",
								X"3F",X"F8",X"38",X"38",X"30",X"18",X"70",X"1C",
								X"70",X"1C",X"60",X"1C",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"C0", -- B
								X"7F",X"F0",X"71",X"F8",X"70",X"38",X"70",X"38",  -- 11
								X"70",X"38",X"70",X"38",X"71",X"F0",X"7F",X"E0",
								X"7F",X"F0",X"70",X"78",X"70",X"3C",X"70",X"1C",
								X"70",X"1C",X"70",X"1C",X"70",X"3C",X"71",X"F8",
								X"7F",X"F0",X"7F",X"C0",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"E0", -- C
								X"0F",X"F8",X"1F",X"7C",X"3C",X"1C",X"38",X"08",  -- 12
								X"38",X"00",X"70",X"00",X"70",X"00",X"70",X"00",
								X"70",X"00",X"70",X"00",X"70",X"00",X"70",X"00",
								X"78",X"00",X"38",X"00",X"3C",X"1C",X"1F",X"7C",
								X"0F",X"F8",X"03",X"E0",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"80", -- D
								X"7F",X"E0",X"71",X"F0",X"70",X"78",X"70",X"38",  -- 13
								X"70",X"1C",X"70",X"1C",X"70",X"1C",X"70",X"1C",
								X"70",X"1C",X"70",X"1C",X"70",X"1C",X"70",X"1C",
								X"70",X"1C",X"70",X"38",X"70",X"78",X"71",X"F0",
								X"7F",X"E0",X"7F",X"80",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"FC", -- E
								X"3F",X"FC",X"30",X"00",X"30",X"00",X"30",X"00",  -- 14
								X"30",X"00",X"30",X"00",X"3F",X"F0",X"3F",X"F0",
								X"3F",X"F0",X"30",X"00",X"30",X"00",X"30",X"00",
								X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",
								X"3F",X"F8",X"3F",X"F8",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"F8", -- F
								X"3F",X"F8",X"38",X"00",X"38",X"00",X"38",X"00",  -- 15
								X"38",X"00",X"38",X"00",X"38",X"00",X"3F",X"F0",
								X"3F",X"F0",X"38",X"00",X"38",X"00",X"38",X"00",
								X"38",X"00",X"38",X"00",X"38",X"00",X"38",X"00",
								X"38",X"00",X"38",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"E0", -- G
								X"0F",X"F8",X"1F",X"FC",X"3C",X"1C",X"38",X"08",  -- 16
								X"70",X"00",X"70",X"00",X"70",X"00",X"70",X"00",
								X"70",X"00",X"70",X"FC",X"70",X"FC",X"70",X"1C",
								X"70",X"1C",X"38",X"1C",X"3C",X"1C",X"1F",X"7C",
								X"0F",X"FC",X"07",X"E0",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"1C", -- H
								X"70",X"1C",X"70",X"1C",X"70",X"1C",X"70",X"1C",  -- 17
								X"70",X"1C",X"70",X"1C",X"70",X"1C",X"7F",X"FC",
								X"7F",X"FC",X"70",X"1C",X"70",X"1C",X"70",X"1C",
								X"70",X"1C",X"70",X"1C",X"70",X"1C",X"70",X"1C",
								X"70",X"1C",X"70",X"1C",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"F0", -- I
								X"3F",X"F0",X"03",X"80",X"03",X"80",X"03",X"80",  -- 18
								X"03",X"80",X"03",X"80",X"03",X"80",X"03",X"80",
								X"03",X"80",X"03",X"80",X"03",X"80",X"03",X"80",
								X"03",X"80",X"03",X"80",X"03",X"80",X"03",X"80",
								X"3F",X"F8",X"3F",X"F8",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"FC", -- J
								X"07",X"FC",X"00",X"E0",X"00",X"E0",X"00",X"E0",  -- 19
								X"00",X"E0",X"00",X"E0",X"00",X"E0",X"00",X"E0",
								X"00",X"E0",X"00",X"E0",X"00",X"E0",X"00",X"E0",
								X"00",X"E0",X"00",X"E0",X"31",X"E0",X"7F",X"C0",
								X"3F",X"80",X"1F",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"70",X"3C",X"70",X"38", -- K
								X"70",X"70",X"70",X"E0",X"71",X"C0",X"73",X"C0",  -- 20
								X"77",X"80",X"77",X"00",X"7F",X"00",X"7F",X"00",
								X"7B",X"80",X"73",X"C0",X"71",X"C0",X"70",X"E0",
								X"70",X"F0",X"70",X"70",X"70",X"78",X"70",X"3C",
								X"70",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"00", -- L
								X"38",X"00",X"38",X"00",X"38",X"00",X"38",X"00",  -- 21
								X"38",X"00",X"38",X"00",X"38",X"00",X"38",X"00",
								X"38",X"00",X"38",X"00",X"38",X"00",X"38",X"00",
								X"38",X"00",X"38",X"00",X"38",X"00",X"38",X"00",
								X"3F",X"FC",X"3F",X"FC",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"70",X"1C",X"70",X"1C", -- M
								X"78",X"3C",X"78",X"3C",X"7C",X"3C",X"7C",X"7C",  -- 22
								X"7C",X"7C",X"76",X"DC",X"76",X"DC",X"77",X"DC",
								X"73",X"9C",X"73",X"9C",X"71",X"1C",X"70",X"1C",
								X"70",X"1C",X"70",X"1C",X"70",X"1C",X"70",X"1C",
								X"70",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"78",X"1C", -- N
								X"78",X"1C",X"7C",X"1C",X"7C",X"1C",X"7E",X"1C",  -- 23
								X"7E",X"1C",X"77",X"1C",X"77",X"1C",X"73",X"9C",
								X"73",X"9C",X"71",X"DC",X"71",X"DC",X"70",X"FC",
								X"70",X"FC",X"70",X"7C",X"70",X"7C",X"70",X"3C",
								X"70",X"3C",X"70",X"1C",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"C0", -- O
								X"1F",X"F0",X"3E",X"F8",X"38",X"38",X"78",X"3C",  -- 24
								X"70",X"1C",X"70",X"1C",X"70",X"1C",X"70",X"1C",
								X"70",X"1C",X"70",X"1C",X"70",X"1C",X"70",X"1C",
								X"70",X"1C",X"70",X"1C",X"38",X"38",X"3E",X"F8",
								X"1F",X"F0",X"07",X"C0",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"E0", -- P
								X"3F",X"F0",X"3F",X"F8",X"38",X"3C",X"38",X"1C",  -- 25
								X"38",X"1C",X"38",X"1C",X"38",X"3C",X"38",X"F8",
								X"3F",X"F0",X"3F",X"E0",X"38",X"00",X"38",X"00",
								X"38",X"00",X"38",X"00",X"38",X"00",X"38",X"00",
								X"38",X"00",X"38",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"C0", -- Q
								X"1F",X"F0",X"1E",X"F8",X"38",X"38",X"78",X"3C",  -- 26
								X"70",X"1C",X"70",X"1C",X"70",X"1C",X"70",X"1C",
								X"70",X"1C",X"70",X"1C",X"70",X"1C",X"70",X"1C",
								X"70",X"1C",X"78",X"1C",X"38",X"38",X"3E",X"F8",
								X"1F",X"F0",X"07",X"C0",X"03",X"80",X"03",X"80",
								X"01",X"E8",X"01",X"F8"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"E0", -- R
								X"7F",X"F0",X"7F",X"F8",X"70",X"38",X"70",X"3C",  -- 27
								X"70",X"1C",X"70",X"1C",X"70",X"38",X"70",X"F8",
								X"7F",X"F0",X"7F",X"E0",X"71",X"C0",X"70",X"E0",
								X"70",X"E0",X"70",X"70",X"70",X"70",X"70",X"38",
								X"70",X"38",X"70",X"1C",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"E0", -- S
								X"1F",X"F0",X"3E",X"F8",X"38",X"10",X"38",X"10",  -- 28
								X"38",X"00",X"3C",X"00",X"1F",X"00",X"0F",X"C0",
								X"07",X"F0",X"01",X"F8",X"00",X"78",X"00",X"1C",
								X"00",X"1C",X"20",X"1C",X"30",X"38",X"7F",X"F8",
								X"3F",X"F0",X"0F",X"C0",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"FC", -- T
								X"7F",X"FC",X"7F",X"FC",X"03",X"80",X"03",X"80",  -- 29
								X"03",X"80",X"03",X"80",X"03",X"80",X"03",X"80",
								X"03",X"80",X"03",X"80",X"03",X"80",X"03",X"80",
								X"03",X"80",X"03",X"80",X"03",X"80",X"03",X"80",
								X"03",X"80",X"03",X"80",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"1C", -- U
								X"70",X"1C",X"70",X"1C",X"70",X"1C",X"70",X"1C",  -- 30
								X"70",X"1C",X"70",X"1C",X"70",X"1C",X"70",X"1C",
								X"70",X"1C",X"70",X"1C",X"70",X"1C",X"70",X"1C",
								X"70",X"1C",X"78",X"1C",X"38",X"38",X"3E",X"F8",
								X"1F",X"F0",X"07",X"C0",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"70",X"0C",X"70",X"1C", -- V
								X"70",X"1C",X"38",X"18",X"38",X"38",X"38",X"38",  -- 31
								X"1C",X"38",X"1C",X"30",X"1C",X"70",X"0C",X"70",
								X"0E",X"60",X"0E",X"E0",X"06",X"E0",X"07",X"C0",
								X"07",X"C0",X"03",X"C0",X"03",X"80",X"03",X"80",
								X"01",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"0E", -- W
								X"61",X"8E",X"61",X"8C",X"63",X"8C",X"73",X"8C",  -- 32
								X"73",X"CC",X"73",X"CC",X"72",X"CC",X"36",X"DC",
								X"36",X"F8",X"36",X"78",X"36",X"78",X"3C",X"78",
								X"3C",X"78",X"3C",X"78",X"1C",X"38",X"18",X"38",
								X"18",X"30",X"18",X"30",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"1C", -- X
								X"38",X"38",X"38",X"38",X"1C",X"70",X"1C",X"70",  -- 33
								X"0E",X"E0",X"0E",X"E0",X"07",X"C0",X"03",X"C0",
								X"03",X"80",X"07",X"C0",X"07",X"C0",X"0E",X"E0",
								X"0E",X"E0",X"1C",X"70",X"1C",X"70",X"38",X"38",
								X"38",X"3C",X"70",X"1C",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"1C", -- Y
								X"70",X"1C",X"38",X"38",X"38",X"38",X"1C",X"70",  -- 34
								X"1C",X"70",X"0E",X"70",X"0E",X"E0",X"07",X"E0",
								X"07",X"C0",X"03",X"C0",X"03",X"80",X"03",X"80",
								X"03",X"80",X"03",X"80",X"03",X"80",X"03",X"80",
								X"03",X"80",X"03",X"80",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"FC", -- Z
								X"3F",X"FC",X"3F",X"F8",X"00",X"38",X"00",X"70",  -- 35
								X"00",X"F0",X"00",X"E0",X"01",X"C0",X"01",X"C0",
								X"03",X"80",X"07",X"80",X"07",X"00",X"0E",X"00",
								X"1E",X"00",X"1C",X"00",X"3C",X"00",X"3F",X"FC",
								X"7F",X"FC",X"7F",X"FC",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- a
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 36
								X"0F",X"C0",X"1F",X"F0",X"3C",X"F8",X"10",X"38",
								X"00",X"38",X"07",X"F8",X"1F",X"F8",X"3C",X"18",
								X"78",X"38",X"70",X"38",X"70",X"38",X"78",X"F8",
								X"3F",X"F8",X"1F",X"B8",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"38",X"00",X"38",X"00", -- b
								X"38",X"00",X"38",X"00",X"38",X"00",X"38",X"00",  -- 37
								X"3B",X"E0",X"3F",X"F0",X"3E",X"F8",X"3C",X"38",
								X"38",X"1C",X"38",X"1C",X"38",X"1C",X"38",X"1C",
								X"38",X"1C",X"38",X"1C",X"38",X"38",X"3E",X"F8",
								X"37",X"F0",X"33",X"E0",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- c
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 38
								X"03",X"E0",X"0F",X"F8",X"1F",X"7C",X"3C",X"18",
								X"38",X"00",X"78",X"00",X"70",X"00",X"70",X"00",
								X"78",X"00",X"38",X"00",X"3C",X"18",X"1F",X"FC",
								X"0F",X"F8",X"03",X"E0",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"3C",X"00",X"38", -- d
								X"00",X"38",X"00",X"38",X"00",X"38",X"00",X"38",  -- 39
								X"07",X"B8",X"1F",X"F8",X"3E",X"F8",X"38",X"38",
								X"70",X"38",X"70",X"38",X"70",X"38",X"70",X"38",
								X"70",X"38",X"78",X"38",X"38",X"38",X"3E",X"F8",
								X"1F",X"F8",X"07",X"9C",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- e
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 40
								X"07",X"C0",X"0F",X"F0",X"1E",X"70",X"38",X"38",
								X"38",X"38",X"70",X"18",X"7F",X"FC",X"7F",X"FC",
								X"70",X"00",X"30",X"00",X"38",X"10",X"1E",X"38",
								X"0F",X"F0",X"07",X"E0",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"01",X"F8",X"03",X"FC", -- f
								X"07",X"9C",X"07",X"04",X"0E",X"00",X"0E",X"00",  -- 41
								X"7F",X"F0",X"7F",X"F0",X"0E",X"00",X"0E",X"00",
								X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",
								X"0E",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00",
								X"0E",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- g
								X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"9C",  -- 42
								X"1F",X"FC",X"3C",X"F0",X"38",X"70",X"30",X"70",
								X"38",X"70",X"3C",X"E0",X"1F",X"E0",X"1F",X"80",
								X"30",X"00",X"38",X"00",X"3F",X"F0",X"1F",X"F8",
								X"30",X"78",X"60",X"1C",X"60",X"1C",X"78",X"78",
								X"3F",X"F0",X"0F",X"C0"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"38",X"00",X"38",X"00", -- h
								X"38",X"00",X"38",X"00",X"38",X"00",X"38",X"00",  -- 43
								X"39",X"E0",X"3B",X"F0",X"3F",X"78",X"3C",X"38",
								X"38",X"38",X"38",X"38",X"38",X"38",X"38",X"38",
								X"38",X"38",X"38",X"38",X"38",X"38",X"38",X"38",
								X"38",X"38",X"38",X"38",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"03",X"00",X"03",X"80", -- i
								X"03",X"80",X"03",X"80",X"00",X"00",X"00",X"00",  -- 44
								X"1F",X"80",X"1F",X"80",X"03",X"80",X"03",X"80",
								X"03",X"80",X"03",X"80",X"03",X"80",X"03",X"80",
								X"03",X"80",X"03",X"80",X"03",X"80",X"03",X"80",
								X"1F",X"F0",X"1F",X"F0",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"40",X"00",X"E0",X"00",X"E0", -- j
								X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",  -- 45
								X"1F",X"E0",X"1F",X"E0",X"00",X"E0",X"00",X"E0",
								X"00",X"E0",X"00",X"E0",X"00",X"E0",X"00",X"E0",
								X"00",X"E0",X"00",X"E0",X"00",X"E0",X"00",X"E0",
								X"00",X"E0",X"00",X"E0",X"00",X"E0",X"30",X"E0",
								X"7F",X"E0",X"3F",X"C0"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"38",X"00",X"38",X"00", -- k
								X"38",X"00",X"38",X"00",X"38",X"00",X"38",X"00",  -- 46
								X"38",X"38",X"38",X"70",X"38",X"E0",X"39",X"C0",
								X"3B",X"80",X"3F",X"00",X"3F",X"80",X"3F",X"C0",
								X"39",X"C0",X"38",X"E0",X"38",X"F0",X"38",X"78",
								X"38",X"38",X"38",X"1C",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"3F",X"80",X"3F",X"80", -- l
								X"03",X"80",X"03",X"80",X"03",X"80",X"03",X"80",  -- 47
								X"03",X"80",X"03",X"80",X"03",X"80",X"03",X"80",
								X"03",X"80",X"03",X"80",X"03",X"80",X"03",X"80",
								X"03",X"80",X"03",X"80",X"03",X"80",X"03",X"80",
								X"3F",X"F8",X"3F",X"F8",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- m
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 48
								X"77",X"38",X"7F",X"7C",X"73",X"DC",X"73",X"8C",
								X"73",X"8C",X"73",X"8C",X"73",X"8C",X"73",X"8C",
								X"73",X"8C",X"73",X"8C",X"73",X"8C",X"73",X"8C",
								X"73",X"8C",X"73",X"8C",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- n
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 49
								X"39",X"E0",X"3B",X"F0",X"3F",X"78",X"3C",X"38",
								X"38",X"38",X"38",X"38",X"38",X"38",X"38",X"38",
								X"38",X"38",X"38",X"38",X"38",X"38",X"38",X"38",
								X"38",X"38",X"38",X"38",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- o
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 50
								X"07",X"C0",X"1F",X"F0",X"3E",X"F8",X"38",X"38",
								X"70",X"1C",X"70",X"1C",X"70",X"1C",X"70",X"1C",
								X"70",X"1C",X"70",X"3C",X"38",X"38",X"3E",X"F8",
								X"1F",X"F0",X"07",X"C0",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- p
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 51
								X"3B",X"E0",X"3F",X"F0",X"3E",X"78",X"38",X"3C",
								X"38",X"1C",X"38",X"1C",X"38",X"1C",X"38",X"1C",
								X"38",X"1C",X"38",X"1C",X"38",X"38",X"3E",X"F8",
								X"3F",X"F0",X"3B",X"E0",X"38",X"00",X"38",X"00",
								X"38",X"00",X"38",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- q
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 52
								X"07",X"9C",X"1F",X"DC",X"3E",X"FC",X"38",X"3C",
								X"70",X"3C",X"70",X"3C",X"70",X"3C",X"70",X"3C",
								X"70",X"3C",X"70",X"3C",X"38",X"3C",X"3E",X"FC",
								X"1F",X"FC",X"0F",X"BC",X"00",X"3C",X"00",X"3C",
								X"00",X"3C",X"00",X"3C"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- r
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 53
								X"1C",X"F0",X"1D",X"FC",X"1F",X"F8",X"1E",X"08",
								X"1C",X"00",X"1C",X"00",X"1C",X"00",X"1C",X"00",
								X"1C",X"00",X"1C",X"00",X"1C",X"00",X"1C",X"00",
								X"1C",X"00",X"1C",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- s
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 54
								X"07",X"E0",X"1F",X"F0",X"3E",X"78",X"38",X"10",
								X"3C",X"00",X"1F",X"00",X"0F",X"E0",X"03",X"F0",
								X"00",X"78",X"00",X"18",X"30",X"18",X"3E",X"78",
								X"3F",X"F0",X"0F",X"E0",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- t
								X"07",X"00",X"07",X"00",X"07",X"00",X"07",X"00",  -- 55
								X"3F",X"F0",X"3F",X"F0",X"07",X"00",X"07",X"00",
								X"07",X"00",X"07",X"00",X"07",X"00",X"07",X"00",
								X"07",X"00",X"07",X"00",X"07",X"08",X"07",X"B8",
								X"03",X"F8",X"01",X"F0",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- u
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 56
								X"38",X"38",X"38",X"38",X"38",X"38",X"38",X"38",
								X"38",X"38",X"38",X"38",X"38",X"38",X"38",X"38",
								X"38",X"38",X"38",X"38",X"38",X"78",X"3C",X"F8",
								X"1F",X"F8",X"0F",X"98",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- v
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 57
								X"70",X"1C",X"38",X"1C",X"38",X"18",X"38",X"38",
								X"1C",X"38",X"1C",X"30",X"1C",X"70",X"0E",X"60",
								X"0E",X"E0",X"07",X"E0",X"07",X"C0",X"07",X"C0",
								X"03",X"80",X"03",X"80",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- w
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 58
								X"E0",X"0E",X"61",X"8C",X"63",X"8C",X"73",X"8C",
								X"73",X"8C",X"73",X"CC",X"32",X"DC",X"36",X"DC",
								X"36",X"F8",X"3E",X"78",X"3C",X"78",X"1C",X"78",
								X"1C",X"78",X"1C",X"30",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- x
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 59
								X"78",X"38",X"38",X"78",X"1C",X"70",X"1E",X"E0",
								X"0E",X"E0",X"07",X"C0",X"03",X"80",X"07",X"C0",
								X"07",X"C0",X"0E",X"E0",X"1E",X"F0",X"1C",X"70",
								X"38",X"38",X"78",X"3C",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- y
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 60
								X"70",X"18",X"38",X"38",X"38",X"38",X"38",X"38",
								X"1C",X"30",X"1C",X"70",X"0E",X"70",X"0E",X"60",
								X"06",X"E0",X"07",X"E0",X"07",X"C0",X"03",X"C0",
								X"03",X"80",X"01",X"80",X"03",X"80",X"03",X"00",
								X"6F",X"00",X"7E",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- z
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  -- 61
								X"3F",X"F8",X"3F",X"F8",X"3F",X"F8",X"00",X"F0",
								X"00",X"E0",X"01",X"C0",X"03",X"80",X"07",X"00",
								X"0F",X"00",X"1E",X"00",X"1C",X"00",X"38",X"0C",
								X"7F",X"FC",X"7F",X"FC",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"03",X"C0",X"03",X"C0",X"03",X"C0", --!
								X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",  --62
								X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",
								X"03",X"C0",X"03",X"C0",X"03",X"C0",X"03",X"C0",
								X"03",X"C0",X"03",X"C0",X"00",X"00",X"00",X"00",
								X"00",X"00",X"03",X"C0",X"03",X"C0",X"03",X"C0",
								X"03",X"C0",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"0C",X"30",X"0C",X"30", --"
								X"0C",X"30",X"0C",X"30",X"0C",X"30",X"0C",X"30",  --63
								X"0C",X"30",X"0C",X"30",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --#
								X"01",X"08",X"03",X"18",X"03",X"18",X"02",X"10",  --64
								X"02",X"10",X"3F",X"FE",X"06",X"30",X"06",X"30",
								X"04",X"20",X"04",X"20",X"04",X"60",X"7F",X"FC",
								X"0C",X"60",X"08",X"40",X"08",X"40",X"18",X"C0",
								X"18",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --%
								X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"10",  --65
								X"44",X"30",X"42",X"20",X"42",X"40",X"42",X"C0",
								X"44",X"80",X"39",X"38",X"03",X"44",X"02",X"42",
								X"04",X"42",X"04",X"42",X"08",X"44",X"10",X"38",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --&
								X"00",X"00",X"00",X"00",X"0F",X"00",X"19",X"80",  --66
								X"10",X"80",X"10",X"88",X"19",X"88",X"0E",X"08",
								X"1B",X"08",X"20",X"88",X"60",X"50",X"60",X"70",
								X"60",X"70",X"30",X"D0",X"1F",X"0E",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --'
								X"01",X"80",X"01",X"80",X"01",X"80",X"01",X"80",  --67
								X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --(
								X"00",X"00",X"00",X"00",X"00",X"C0",X"01",X"80",  --68
								X"01",X"00",X"01",X"00",X"03",X"00",X"02",X"00",
								X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",
								X"02",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
								X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --)
								X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"80",  --69
								X"00",X"80",X"00",X"40",X"00",X"40",X"00",X"40",
								X"00",X"40",X"00",X"40",X"00",X"40",X"00",X"40",
								X"00",X"40",X"00",X"40",X"00",X"80",X"00",X"80",
								X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --*
								X"00",X"80",X"00",X"00",X"06",X"20",X"01",X"80",  --70
								X"02",X"40",X"02",X"40",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --+
								X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"80",  --71
								X"01",X"80",X"01",X"80",X"01",X"80",X"1F",X"F8",
								X"1F",X"F8",X"01",X"80",X"01",X"80",X"01",X"80",
								X"01",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --,
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  --72
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"C0",X"01",X"C0",
								X"01",X"80",X"03",X"00",X"03",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- -
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  --73
								X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"E0",
								X"07",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --.
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  --74
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"03",X"80",X"03",X"80",X"03",X"80",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18", --/
								X"00",X"30",X"00",X"30",X"00",X"20",X"00",X"60",  --75
								X"00",X"60",X"00",X"C0",X"00",X"C0",X"00",X"80",
								X"01",X"80",X"01",X"80",X"03",X"00",X"03",X"00",
								X"02",X"00",X"06",X"00",X"04",X"00",X"0C",X"00",
								X"0C",X"00",X"08",X"00",X"18",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --:
								X"00",X"00",X"00",X"00",X"03",X"80",X"03",X"80",  --76
								X"03",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"80",
								X"03",X"80",X"03",X"80",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --;
								X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",  --77
								X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
								X"00",X"80",X"01",X"80",X"01",X"00",X"01",X"00",
								X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --<
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  --78
								X"00",X"00",X"00",X"30",X"00",X"E0",X"01",X"C0",
								X"07",X"00",X"1C",X"00",X"1C",X"00",X"07",X"00",
								X"01",X"C0",X"00",X"30",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --=
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  --79
								X"00",X"00",X"00",X"00",X"1F",X"FC",X"1F",X"F8",
								X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"FC",
								X"1F",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -->
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  --80
								X"08",X"00",X"0E",X"00",X"03",X"80",X"00",X"E0",
								X"00",X"38",X"00",X"38",X"00",X"70",X"01",X"C0",
								X"07",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --?
								X"01",X"80",X"07",X"E0",X"0E",X"F0",X"00",X"30",  --81
								X"00",X"10",X"00",X"30",X"00",X"20",X"00",X"40",
								X"00",X"80",X"01",X"80",X"01",X"00",X"01",X"00",
								X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"80",
								X"01",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --*C
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",  --82
								X"3C",X"00",X"24",X"00",X"24",X"00",X"24",X"00",
								X"3C",X"00",X"00",X"FC",X"00",X"80",X"00",X"80",
								X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",
								X"00",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --delta
								X"10",X"00",X"18",X"00",X"1C",X"00",X"1E",X"00",  --83
								X"1F",X"00",X"1F",X"80",X"1F",X"C0",X"1F",X"E0",
								X"1F",X"F0",X"1F",X"F8",X"1F",X"F0",X"1F",X"E0",
								X"1F",X"C0",X"1F",X"00",X"1E",X"00",X"18",X"00",
								X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --||
								X"00",X"00",X"00",X"00",X"0E",X"38",X"0E",X"38",  --84
								X"0E",X"38",X"0E",X"38",X"0E",X"38",X"0E",X"38",
								X"0E",X"38",X"0E",X"38",X"0E",X"38",X"0E",X"38",
								X"0E",X"38",X"0E",X"38",X"0E",X"38",X"0E",X"38",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								X"00",X"00",X"00",X"00")
								);
    --------------------------------------------------------------------------------
	-- 0~9 A~Z a~z
	type rom16x12 is array (0 to 84, 0 to 31) of std_logic_vector(7 downto 0); -- rows x cols
	constant Font16 : rom16x12 :=( -- 16 x 16 / 8 = 32 Bytes (Padding to 16 x 16)
								-------------------------------------------------
								(X"00",X"00",X"0E",X"00",X"1B",X"00",X"31",X"80", -- 0
								 X"31",X"80",X"33",X"80",X"26",X"80",X"24",X"80", -- 0
								 X"39",X"80",X"31",X"80",X"31",X"80",X"1B",X"00",
								 X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"0E",X"00",X"1E",X"00",X"06",X"00", -- 1
								 X"06",X"00",X"06",X"00",X"06",X"00",X"06",X"00", -- 1
								 X"06",X"00",X"06",X"00",X"06",X"00",X"06",X"00",
								 X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"1E",X"00",X"3F",X"00",X"31",X"80", -- 2
								 X"01",X"80",X"01",X"80",X"01",X"80",X"03",X"00", -- 2
								 X"06",X"00",X"0C",X"00",X"18",X"00",X"30",X"00",
								 X"3F",X"80",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"1E",X"00",X"3B",X"00",X"01",X"80", -- 3
								 X"01",X"00",X"07",X"00",X"0E",X"00",X"03",X"00", -- 3
								 X"01",X"80",X"01",X"80",X"01",X"80",X"3B",X"00",
								 X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"03",X"00",X"03",X"00",X"07",X"00", -- 4
								 X"0F",X"00",X"0B",X"00",X"1B",X"00",X"13",X"00", -- 4
								 X"33",X"00",X"3F",X"C0",X"03",X"00",X"03",X"00",
								 X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"1F",X"80",X"10",X"00",X"10",X"00", -- 5
								 X"10",X"00",X"1F",X"00",X"3B",X"80",X"01",X"80", -- 5
								 X"01",X"80",X"01",X"80",X"11",X"80",X"3B",X"00",
								 X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"0F",X"00",X"1F",X"00",X"10",X"00", -- 6
								 X"30",X"00",X"3F",X"00",X"3B",X"80",X"31",X"80", -- 6
								 X"31",X"80",X"31",X"80",X"31",X"80",X"1B",X"00",
								 X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"3F",X"80",X"3F",X"80",X"01",X"00", -- 7
								 X"03",X"00",X"03",X"00",X"06",X"00",X"06",X"00", -- 7
								 X"06",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",
								 X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"0F",X"00",X"1B",X"00",X"31",X"80", -- 8
								 X"31",X"80",X"1B",X"00",X"0E",X"00",X"1B",X"00", -- 8
								 X"31",X"80",X"31",X"80",X"31",X"80",X"3F",X"80",
								 X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"0E",X"00",X"1B",X"00",X"31",X"80", -- 9
								X"31",X"80",X"31",X"80",X"31",X"80",X"1B",X"80",  -- 9
								X"0F",X"80",X"01",X"80",X"01",X"00",X"3F",X"00",
								X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"04",X"00",X"04",X"00",X"0E",X"00", -- A
								 X"0E",X"00",X"0A",X"00",X"1B",X"00",X"1B",X"00", -- 10
								 X"11",X"00",X"3F",X"80",X"31",X"80",X"20",X"80",
								 X"60",X"C0",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"3F",X"00",X"33",X"80",X"31",X"80", -- B
								 X"31",X"80",X"33",X"00",X"3F",X"00",X"31",X"80", -- 11
								 X"31",X"80",X"30",X"80",X"31",X"80",X"3F",X"80",
								 X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"0F",X"00",X"1D",X"80",X"30",X"80", -- C
								X"30",X"00",X"20",X"00",X"20",X"00",X"20",X"00",  -- 12
								X"20",X"00",X"30",X"00",X"30",X"80",X"1F",X"80",
								X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"3E",X"00",X"37",X"00",X"31",X"80", -- D
								 X"31",X"80",X"30",X"80",X"30",X"80",X"30",X"80", -- 13
								 X"30",X"80",X"31",X"80",X"31",X"80",X"37",X"00",
								 X"3E",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"3F",X"80",X"30",X"00",X"30",X"00", -- E
								 X"30",X"00",X"30",X"00",X"3F",X"00",X"3F",X"00", -- 14
								 X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",
								 X"3F",X"80",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"3F",X"80",X"30",X"00",X"30",X"00", -- F
								 X"30",X"00",X"30",X"00",X"3F",X"00",X"30",X"00", -- 15
								 X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",
								 X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"0F",X"00",X"1F",X"80",X"30",X"80", -- G
								 X"30",X"00",X"20",X"00",X"20",X"00",X"23",X"80", -- 16
								 X"20",X"80",X"30",X"80",X"30",X"80",X"1F",X"80",
								 X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"31",X"80",X"31",X"80",X"31",X"80", -- H
								 X"31",X"80",X"31",X"80",X"3F",X"80",X"31",X"80", -- 17
								 X"31",X"80",X"31",X"80",X"31",X"80",X"31",X"80",
								 X"31",X"80",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"3F",X"00",X"04",X"00",X"04",X"00", -- I
								 X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00", -- 18
								 X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",
								 X"3F",X"80",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"0F",X"80",X"03",X"00",X"03",X"00", -- J
								 X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00", -- 19
								 X"03",X"00",X"03",X"00",X"02",X"00",X"3E",X"00",
								 X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"21",X"80",X"23",X"00",X"23",X"00",X"26",X"00", -- K
								X"2C",X"00",X"3C",X"00",X"3C",X"00",X"26",X"00",  -- 20
								X"23",X"00",X"23",X"00",X"21",X"80",X"21",X"80",
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"30",X"00",X"30",X"00",X"30",X"00", -- L
								 X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00", -- 21
								 X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",
								 X"3F",X"80",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"20",X"80",X"31",X"80",X"31",X"80",X"3B",X"80", -- M
								 X"2A",X"80",X"2A",X"80",X"2E",X"80",X"24",X"80", -- 22
								 X"20",X"80",X"20",X"80",X"20",X"80",X"20",X"80",
								 X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"30",X"80",X"30",X"80",X"38",X"80", -- N
								X"38",X"80",X"2C",X"80",X"2C",X"80",X"26",X"80",  -- 23
								X"26",X"80",X"23",X"80",X"23",X"80",X"21",X"80",
								X"21",X"80",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"0E",X"00",X"3B",X"80",X"31",X"80", -- O
								X"20",X"80",X"60",X"C0",X"60",X"C0",X"60",X"C0",  -- 24
								X"60",X"C0",X"20",X"80",X"31",X"80",X"3B",X"80",
								X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"3F",X"00",X"3F",X"80",X"31",X"80", -- P
								 X"30",X"80",X"31",X"80",X"3F",X"80",X"3F",X"00", -- 25
								 X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00",
								 X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"0E",X"00",X"1B",X"00",X"31",X"80", -- Q
								 X"20",X"80",X"60",X"C0",X"60",X"C0",X"60",X"C0", -- 26
								 X"60",X"C0",X"20",X"80",X"31",X"80",X"1B",X"80",
								 X"0F",X"00",X"04",X"00",X"06",X"80",X"03",X"80"),
								-------------------------------------------------
								(X"00",X"00",X"3F",X"00",X"3F",X"80",X"31",X"80", -- R
								 X"31",X"80",X"31",X"80",X"3F",X"80",X"3F",X"00", -- 27
								 X"32",X"00",X"33",X"00",X"33",X"00",X"31",X"80",
								 X"31",X"80",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"0F",X"00",X"1B",X"80",X"30",X"00", -- S
								 X"30",X"00",X"38",X"00",X"1E",X"00",X"07",X"80", -- 28
								 X"01",X"80",X"00",X"80",X"21",X"80",X"3F",X"80",
								 X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"7F",X"80",X"7F",X"80",X"04",X"00", -- T
								 X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00", -- 29
								 X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",
								 X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"30",X"80",X"30",X"80",X"30",X"80", -- U
								 X"30",X"80",X"30",X"80",X"30",X"80",X"30",X"80", -- 30
								 X"30",X"80",X"30",X"80",X"31",X"80",X"3B",X"80",
								 X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"20",X"C0",X"30",X"80",X"31",X"80",X"31",X"80", -- V
								 X"11",X"00",X"19",X"00",X"1B",X"00",X"0A",X"00", -- 31
								 X"0E",X"00",X"0E",X"00",X"06",X"00",X"04",X"00",
								 X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"60",X"C0",X"64",X"C0",X"24",X"C0", -- W
								 X"26",X"80",X"2E",X"80",X"2A",X"80",X"3A",X"80", -- 32
								 X"3B",X"80",X"39",X"80",X"31",X"80",X"11",X"80",
								 X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"31",X"80",X"31",X"80",X"1B",X"00", -- X
								 X"1B",X"00",X"0E",X"00",X"0E",X"00",X"0E",X"00", -- 33
								 X"0E",X"00",X"1B",X"00",X"1B",X"00",X"31",X"80",
								 X"31",X"80",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"20",X"80",X"31",X"80",X"11",X"80", -- Y
								 X"1B",X"00",X"1B",X"00",X"0E",X"00",X"0E",X"00", -- 34
								 X"06",X"00",X"06",X"00",X"06",X"00",X"06",X"00",
								 X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"3F",X"80",X"3F",X"80",X"01",X"00", -- Z
								 X"03",X"00",X"06",X"00",X"06",X"00",X"0C",X"00", -- 35
								 X"0C",X"00",X"18",X"00",X"18",X"00",X"3F",X"C0",
								 X"3F",X"C0",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- a
								 X"1F",X"00",X"3B",X"80",X"01",X"80",X"01",X"80", -- 36
								 X"1F",X"80",X"31",X"80",X"31",X"80",X"33",X"80",
								 X"1F",X"80",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00", -- b
								 X"37",X"00",X"3B",X"80",X"31",X"80",X"30",X"80", -- 37
								 X"30",X"80",X"30",X"80",X"31",X"80",X"3B",X"80",
								 X"2F",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- c
								 X"0F",X"00",X"1D",X"80",X"30",X"00",X"30",X"00", -- 38
								 X"30",X"00",X"30",X"00",X"30",X"00",X"1F",X"80",
								 X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"01",X"80",X"01",X"80",X"01",X"80",X"01",X"80", -- d
								 X"1F",X"80",X"3B",X"80",X"31",X"80",X"21",X"80", -- 39
								 X"21",X"80",X"31",X"80",X"31",X"80",X"3B",X"80",
								 X"1F",X"80",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- e
								 X"0E",X"00",X"1B",X"00",X"31",X"80",X"31",X"80", -- 40
								 X"3F",X"80",X"20",X"00",X"30",X"00",X"19",X"80",
								 X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"07",X"80",X"0C",X"80",X"0C",X"00",X"08",X"00", -- f
								 X"3F",X"00",X"08",X"00",X"08",X"00",X"08",X"00", -- 41
								 X"08",X"00",X"08",X"00",X"08",X"00",X"08",X"00",
								 X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"C0", -- g
								 X"3B",X"00",X"31",X"00",X"31",X"00",X"33",X"00", -- 42
								 X"1E",X"00",X"30",X"00",X"3F",X"00",X"3F",X"80",
								 X"20",X"80",X"31",X"80",X"1F",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00", -- h
								 X"37",X"00",X"3B",X"80",X"31",X"80",X"31",X"80", -- 43
								 X"31",X"80",X"31",X"80",X"31",X"80",X"31",X"80",
								 X"31",X"80",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"0E",X"00",X"04",X"00",X"00",X"00",X"1C",X"00", -- i
								 X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00", -- 44
								 X"04",X"00",X"04",X"00",X"04",X"00",X"1F",X"00",
								 X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"03",X"00",X"03",X"00",X"00",X"00",X"00",X"00", -- j
								 X"1F",X"00",X"03",X"00",X"03",X"00",X"03",X"00", -- 45
								 X"03",X"00",X"03",X"00",X"03",X"00",X"03",X"00",
								 X"03",X"00",X"03",X"00",X"3E",X"00",X"1C",X"00"),
								-------------------------------------------------
								(X"30",X"00",X"30",X"00",X"30",X"00",X"30",X"00", -- k
								 X"31",X"80",X"33",X"00",X"36",X"00",X"3C",X"00", -- 46
								 X"3E",X"00",X"36",X"00",X"33",X"00",X"31",X"80",
								 X"31",X"80",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"3C",X"00",X"04",X"00",X"04",X"00",X"04",X"00", -- l
								 X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00", -- 47
								 X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00",
								 X"3F",X"80",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- m
								 X"3D",X"80",X"36",X"80",X"24",X"C0",X"24",X"C0", -- 48
								 X"24",X"C0",X"24",X"C0",X"24",X"C0",X"24",X"C0",
								 X"24",X"C0",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- n
								 X"37",X"00",X"3B",X"80",X"31",X"80",X"31",X"80", -- 49
								 X"31",X"80",X"31",X"80",X"31",X"80",X"31",X"80",
								 X"31",X"80",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- o
								 X"0E",X"00",X"1B",X"00",X"31",X"80",X"20",X"80", -- 50
								 X"20",X"80",X"20",X"80",X"31",X"80",X"3B",X"00",
								 X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- p
								 X"3F",X"00",X"3B",X"80",X"31",X"80",X"30",X"80", -- 51
								 X"30",X"80",X"30",X"80",X"31",X"80",X"3B",X"80",
								 X"3F",X"00",X"30",X"00",X"30",X"00",X"30",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- q
								 X"1F",X"80",X"3B",X"80",X"31",X"80",X"21",X"80", -- 52
								 X"21",X"80",X"21",X"80",X"31",X"80",X"3B",X"80",
								 X"1F",X"80",X"01",X"80",X"01",X"80",X"01",X"80"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- r
								 X"1B",X"80",X"1F",X"80",X"18",X"80",X"18",X"00", -- 53
								 X"18",X"00",X"18",X"00",X"18",X"00",X"18",X"00",
								 X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- s
								 X"1F",X"00",X"1B",X"80",X"30",X"00",X"1C",X"00", -- 54
								 X"0F",X"00",X"01",X"80",X"21",X"80",X"3B",X"80",
								 X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"0C",X"00",X"0C",X"00", -- t
								 X"3F",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00", -- 55
								 X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0D",X"80",
								 X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- u
								 X"31",X"80",X"31",X"80",X"31",X"80",X"31",X"80", -- 56
								 X"31",X"80",X"31",X"80",X"31",X"80",X"3B",X"80",
								 X"1F",X"80",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- v
								 X"30",X"80",X"31",X"80",X"31",X"80",X"19",X"00", -- 57
								 X"1B",X"00",X"0B",X"00",X"0E",X"00",X"0E",X"00",
								 X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- w
								 X"60",X"C0",X"64",X"C0",X"24",X"80",X"26",X"80", -- 58
								 X"2A",X"80",X"3A",X"80",X"3B",X"80",X"1B",X"80",
								 X"11",X"80",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- x
								 X"31",X"80",X"1B",X"00",X"1B",X"00",X"0E",X"00", -- 59
								 X"06",X"00",X"0E",X"00",X"1B",X"00",X"11",X"00",
								 X"31",X"80",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- y
								 X"31",X"80",X"31",X"80",X"11",X"80",X"19",X"00", -- 60
								 X"1B",X"00",X"0A",X"00",X"0E",X"00",X"06",X"00",
								 X"04",X"00",X"04",X"00",X"2C",X"00",X"38",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- z
								 X"3F",X"80",X"3F",X"80",X"03",X"00",X"06",X"00", -- 61
								 X"0C",X"00",X"0C",X"00",X"18",X"00",X"3F",X"80",
								 X"3F",X"80",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"04",X"00",X"04",X"00", --!
								 X"04",X"00",X"04",X"00",X"04",X"00",X"04",X"00", --62
								 X"04",X"00",X"04",X"00",X"04",X"00",X"00",X"00",
								 X"00",X"00",X"04",X"00",X"04",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"09",X"00",X"09",X"00", --"
								 X"09",X"00",X"09",X"00",X"00",X"00",X"00",X"00", --63
								 X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								 X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"80", --#
								 X"08",X"00",X"08",X"00",X"7F",X"E0",X"09",X"00", --64
								 X"01",X"00",X"7F",X"C0",X"12",X"00",X"02",X"00",
								 X"02",X"00",X"22",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"38",X"40",X"48",X"80", --%
								 X"40",X"00",X"49",X"00",X"32",X"00",X"02",X"00", --65
								 X"04",X"E0",X"09",X"00",X"09",X"10",X"11",X"00",
								 X"20",X"E0",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"1C",X"00",X"12",X"00", --&
								 X"22",X"00",X"22",X"00",X"1C",X"00",X"34",X"40", --66
								 X"22",X"40",X"41",X"C0",X"41",X"80",X"41",X"80",
								 X"3E",X"60",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"04",X"00",X"04",X"00",X"04",X"00", --'
								 X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --67
								 X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								 X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"02",X"00",X"00",X"00",X"04",X"00", --(
								 X"00",X"00",X"08",X"00",X"08",X"00",X"08",X"00", --68
								 X"08",X"00",X"08",X"00",X"00",X"00",X"04",X"00",
								 X"04",X"00",X"02",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"04",X"00",X"02",X"00", --)
								 X"02",X"00",X"02",X"00",X"00",X"00",X"00",X"00", --69
								 X"00",X"00",X"00",X"00",X"02",X"00",X"02",X"00",
								 X"02",X"00",X"04",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --*
								 X"0E",X"00",X"06",X"00",X"04",X"00",X"00",X"00", --70
								 X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								 X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --+
								 X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"80", --71
								 X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								 X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --,
								 X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --72
								 X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",
								 X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- -
								 X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00", --73
								 X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								 X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --.
								 X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --74
								 X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								 X"06",X"00",X"06",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"80", --/
								 X"01",X"00",X"01",X"00",X"02",X"00",X"02",X"00", --75
								 X"04",X"00",X"04",X"00",X"04",X"00",X"08",X"00",
								 X"08",X"00",X"10",X"00",X"10",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --:
								 X"02",X"00",X"06",X"00",X"00",X"00",X"00",X"00", --76
								 X"00",X"00",X"00",X"00",X"02",X"00",X"02",X"00",
								 X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00", --;
								 X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --77
								 X"00",X"00",X"04",X"00",X"04",X"00",X"04",X"00",
								 X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --<
								 X"00",X"00",X"01",X"00",X"06",X"00",X"18",X"00", --78
								 X"18",X"00",X"02",X"00",X"00",X"00",X"00",X"00",
								 X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --=
								 X"00",X"00",X"1F",X"80",X"00",X"00",X"00",X"00", --79
								 X"1F",X"80",X"00",X"00",X"00",X"00",X"00",X"00",
								 X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -->
								 X"00",X"00",X"10",X"00",X"0C",X"00",X"03",X"00", --80
								 X"00",X"80",X"03",X"00",X"0C",X"00",X"10",X"00",
								 X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00", --?
								 X"01",X"00",X"01",X"00",X"01",X"00",X"02",X"00", --81
								 X"04",X"00",X"04",X"00",X"00",X"00",X"00",X"00",
								 X"04",X"00",X"04",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- Space
								 X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- 82
								 X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								 X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								-------------------------------------------------
								(X"FF",X"F0",X"FF",X"F0",X"7F",X"E0",X"7F",X"E0", -- Inverted
								 X"3F",X"C0",X"3F",X"C0",X"1F",X"80",X"1F",X"80", -- Triangle
								 X"0F",X"00",X"0F",X"00",X"06",X"00",X"06",X"00", -- 83
								 X"06",X"00",X"06",X"00",X"00",X"00",X"0F",X"00"),
								-------------------------------------------------
								(X"FF",X"F0",X"FF",X"F0",X"FF",X"F0",X"FF",X"F0", -- Square
								 X"FF",X"F0",X"FF",X"F0",X"FF",X"F0",X"FF",X"F0", -- 84
								 X"FF",X"F0",X"FF",X"F0",X"FF",X"F0",X"FF",X"F0",
								 X"FF",X"F0",X"FF",X"F0",X"FF",X"F0",X"FF",X"F0")
								-------------------------------------------------
								);
    --------------------------------------------------------------------------------
	type rom32x16 is array (0 to 15, 0 to 63) of std_logic_vector(7 downto 0); 
	constant Font32 : rom32x16 :=( -- 32 x 16 / 8 = 64 Bytes (rows x cols = H x W)
								----------------------------------------------------
								(X"00",X"00",X"00",X"00", -- Mon
								 X"00",X"00",X"00",X"00", -- 0
								 X"00",X"00",X"00",X"00",
								 X"1C",X"38",X"00",X"00",
								 X"1C",X"78",X"00",X"00",
								 X"1C",X"78",X"C1",X"80",
								 X"3C",X"FB",X"F1",X"F0",
								 X"34",X"B3",X"33",X"F8",
								 X"35",X"B6",X"13",X"18",
								 X"35",X"B6",X"1B",X"18",
								 X"37",X"36",X"1B",X"18",
								 X"77",X"76",X"33",X"38",
								 X"66",X"63",X"F6",X"33",
								 X"66",X"61",X"C6",X"33",
								 X"00",X"00",X"00",X"00",
								 X"00",X"00",X"00",X"00"),
								----------------------------------------------------
								(X"00",X"00",X"00",X"00", -- Tue
								 X"00",X"00",X"00",X"00", -- 1
								 X"1F",X"F8",X"00",X"00",
								 X"3F",X"F0",X"00",X"00",
								 X"03",X"80",X"00",X"00",
								 X"03",X"80",X"00",X"00",
								 X"03",X"80",X"00",X"00",
								 X"03",X"00",X"01",X"C0",
								 X"07",X"06",X"33",X"60",
								 X"07",X"06",X"36",X"30",
								 X"07",X"06",X"37",X"F0",
								 X"0E",X"06",X"37",X"E0",
								 X"0E",X"06",X"36",X"00",
								 X"0E",X"07",X"F3",X"F3",
								 X"0C",X"03",X"E1",X"E3",
								 X"00",X"00",X"00",X"00"),
								----------------------------------------------------
								(X"00",X"00",X"00",X"00", -- Wed
								 X"00",X"00",X"00",X"00", -- 2
								 X"70",X"0C",X"00",X"00",
								 X"73",X"0C",X"00",X"0C",
								 X"33",X"98",X"00",X"0C",
								 X"33",X"98",X"00",X"18",
								 X"33",X"98",X"00",X"18",
								 X"37",X"99",X"C1",X"D8",
								 X"36",X"D3",X"63",X"F8",
								 X"1E",X"F6",X"33",X"38",
								 X"1C",X"F7",X"F6",X"18",
								 X"1C",X"E7",X"F6",X"18",
								 X"0C",X"66",X"06",X"38",
								 X"0C",X"63",X"F3",X"F3",
								 X"00",X"01",X"E1",X"C3",
								 X"00",X"00",X"00",X"00"),
								----------------------------------------------------
								(X"00",X"00",X"00",X"00", -- Thu
								 X"00",X"00",X"00",X"00", -- 3
								 X"3F",X"E6",X"00",X"00",
								 X"7F",X"C6",X"00",X"00",
								 X"06",X"0C",X"00",X"00",
								 X"06",X"0C",X"00",X"00",
								 X"06",X"18",X"00",X"00",
								 X"0C",X"18",X"00",X"00",
								 X"1C",X"1B",X"83",X"18",
								 X"1C",X"1F",X"C7",X"38",
								 X"1C",X"1C",X"C6",X"30",
								 X"1C",X"38",X"C6",X"30",
								 X"18",X"30",X"C6",X"30",
								 X"38",X"31",X"87",X"F3",
								 X"38",X"31",X"83",X"E3",
								 X"00",X"00",X"00",X"00"),
								----------------------------------------------------
								(X"00",X"00",X"00",X"00", -- Fri
								 X"00",X"00",X"00",X"00", -- 4
								 X"1F",X"C0",X"00",X"00",
								 X"1F",X"C0",X"00",X"00",
								 X"1C",X"00",X"00",X"00",
								 X"1C",X"00",X"01",X"80",
								 X"1C",X"0C",X"E1",X"80",
								 X"3F",X"8D",X"E0",X"00",
								 X"3F",X"8F",X"81",X"80",
								 X"38",X"0E",X"01",X"80",
								 X"38",X"0C",X"01",X"80",
								 X"30",X"0C",X"01",X"80",
								 X"30",X"0C",X"01",X"80",
								 X"70",X"0C",X"01",X"83",
								 X"70",X"0C",X"01",X"83",
								 X"00",X"00",X"00",X"00"),
								----------------------------------------------------
								(X"00",X"00",X"00",X"00", -- Sat
								 X"0F",X"00",X"00",X"00", -- 5
								 X"1F",X"80",X"00",X"00",
								 X"39",X"C0",X"01",X"80",
								 X"38",X"C0",X"01",X"80",
								 X"38",X"00",X"01",X"80",
								 X"3C",X"07",X"87",X"F0",
								 X"1E",X"0F",X"87",X"F0",
								 X"07",X"9C",X"C1",X"80",
								 X"03",X"98",X"C1",X"80",
								 X"71",X"D8",X"C1",X"80",
								 X"71",X"D8",X"C1",X"80",
								 X"3F",X"9F",X"C1",X"B0",
								 X"1F",X"0F",X"61",X"F3",
								 X"0E",X"06",X"60",X"E3",
								 X"00",X"00",X"00",X"00"),
								----------------------------------------------------
								(X"00",X"00",X"00",X"00", -- Sun
								 X"0F",X"00",X"00",X"00", -- 6
								 X"1F",X"80",X"00",X"00",
								 X"39",X"C0",X"00",X"00",
								 X"38",X"C0",X"00",X"00",
								 X"38",X"00",X"06",X"00",
								 X"3C",X"0C",X"66",X"60",
								 X"1E",X"1C",X"66",X"F0",
								 X"07",X"98",X"67",X"F0",
								 X"03",X"98",X"67",X"98",
								 X"71",X"D8",X"67",X"18",
								 X"71",X"DC",X"E6",X"18",
								 X"3F",X"8F",X"E6",X"18",
								 X"1F",X"0F",X"6E",X"33",
								 X"0E",X"06",X"6C",X"33",
								 X"00",X"00",X"00",X"00"),
								----------------------------------------------------
								(X"00",X"00",X"00",X"00", -- deg C
								 X"01",X"80",X"00",X"00", -- 7
								 X"02",X"40",X"00",X"00",
								 X"02",X"4F",X"C0",X"00",
								 X"01",X"9F",X"E0",X"00",
								 X"00",X"18",X"60",X"00",
								 X"00",X"30",X"00",X"00",
								 X"00",X"30",X"00",X"00",
								 X"00",X"30",X"00",X"00",
								 X"00",X"30",X"00",X"00",
								 X"00",X"30",X"00",X"00",
								 X"00",X"18",X"60",X"00",
								 X"00",X"1F",X"E0",X"00",
								 X"00",X"07",X"C0",X"00",
								 X"00",X"00",X"00",X"00",
								 X"00",X"00",X"00",X"00"),
								----------------------------------------------------
								(X"00",X"00",X"00",X"00", -- deg F
								 X"01",X"80",X"00",X"00", -- 8
								 X"02",X"40",X"00",X"00",
								 X"02",X"4F",X"E0",X"00",
								 X"01",X"8F",X"E0",X"00",
								 X"00",X"0C",X"00",X"00",
								 X"00",X"0C",X"00",X"00",
								 X"00",X"1C",X"00",X"00",
								 X"00",X"1F",X"C0",X"00",
								 X"00",X"1F",X"C0",X"00",
								 X"00",X"1C",X"00",X"00",
								 X"00",X"1C",X"00",X"00",
								 X"00",X"38",X"00",X"00",
								 X"00",X"38",X"00",X"00",
								 X"00",X"38",X"00",X"00",
								 X"00",X"00",X"00",X"00"),
								----------------------------------------------------
								(X"00",X"00",X"00",X"00", -- RH
								 X"00",X"00",X"00",X"00", -- 9
								 X"01",X"F8",X"18",X"30",
								 X"03",X"FC",X"18",X"30",
								 X"03",X"9C",X"18",X"30",
								 X"07",X"1C",X"38",X"70",
								 X"07",X"38",X"30",X"60",
								 X"0F",X"F0",X"30",X"60",
								 X"0F",X"C0",X"7F",X"E0",
								 X"0F",X"C0",X"7F",X"E0",
								 X"0C",X"E0",X"60",X"C0",
								 X"1C",X"70",X"60",X"C0",
								 X"1C",X"30",X"E1",X"C0",
								 X"18",X"30",X"E1",X"C0",
								 X"00",X"00",X"C1",X"80",
								 X"00",X"00",X"00",X"00"),
								----------------------------------------------------
								(X"00",X"00",X"00",X"00", -- percent(%)
								 X"00",X"70",X"0C",X"00", -- 10
								 X"00",X"88",X"1C",X"00",
								 X"00",X"88",X"38",X"00",
								 X"00",X"88",X"70",X"00",
								 X"00",X"70",X"E0",X"00",
								 X"00",X"01",X"C0",X"00",
								 X"00",X"03",X"80",X"00",
								 X"00",X"07",X"00",X"00",
								 X"00",X"0E",X"00",X"00",
								 X"00",X"1C",X"38",X"00",
								 X"00",X"38",X"44",X"00",
								 X"00",X"70",X"44",X"00",
								 X"00",X"E0",X"44",X"00",
								 X"00",X"C0",X"38",X"00",
								 X"00",X"00",X"00",X"00"),
								----------------------------------------------------
								(X"00",X"00",X"00",X"00", -- colon(:)
								 X"00",X"00",X"00",X"00", -- 11
								 X"00",X"01",X"80",X"00",
								 X"00",X"03",X"C0",X"00",
								 X"00",X"03",X"C0",X"00",
								 X"00",X"01",X"80",X"00",
								 X"00",X"00",X"00",X"00",
								 X"00",X"00",X"00",X"00",
								 X"00",X"00",X"00",X"00",
								 X"00",X"00",X"00",X"00",
								 X"00",X"01",X"80",X"00",
								 X"00",X"03",X"C0",X"00",
								 X"00",X"03",X"C0",X"00",
								 X"00",X"01",X"80",X"00",
								 X"00",X"00",X"00",X"00",
								 X"00",X"00",X"00",X"00"),
								----------------------------------------------------
								(X"00",X"00",X"00",X"00", -- ~
								 X"00",X"00",X"00",X"00", -- 12
								 X"00",X"00",X"00",X"00",
								 X"00",X"00",X"00",X"00",
								 X"00",X"00",X"00",X"00",
								 X"00",X"1C",X"00",X"00",
								 X"00",X"3F",X"00",X"00",
								 X"00",X"73",X"80",X"00",
								 X"00",X"C1",X"C1",X"80",
								 X"00",X"00",X"E7",X"00",
								 X"00",X"00",X"7E",X"00",
								 X"00",X"00",X"1C",X"00",
								 X"00",X"00",X"00",X"00",
								 X"00",X"00",X"00",X"00",
								 X"00",X"00",X"00",X"00",
								 X"00",X"00",X"00",X"00"),
								----------------------------------------------------
								(X"00",X"00",X"00",X"00", --vol.
								 X"00",X"00",X"00",X"00", --13
								 X"00",X"00",X"00",X"00",
								 X"04",X"20",X"08",X"00",
								 X"04",X"20",X"04",X"00",
								 X"04",X"20",X"04",X"00",
								 X"04",X"60",X"04",X"00",
								 X"04",X"40",X"04",X"00",
								 X"04",X"CF",X"C4",X"00",
								 X"02",X"8A",X"44",X"00",
								 X"03",X"88",X"44",X"60",
								 X"03",X"08",X"44",X"E0",
								 X"01",X"0E",X"44",X"E0",
								 X"00",X"03",X"80",X"00",
								 X"00",X"00",X"00",X"00",
								 X"00",X"00",X"00",X"00"),
								----------------------------------------------------
								(X"00",X"00",X"00",X"00", --on
								 X"00",X"00",X"00",X"00", --14
								 X"03",X"E0",X"00",X"00",
								 X"02",X"30",X"00",X"00",
								 X"06",X"18",X"00",X"00",
								 X"04",X"08",X"00",X"00",
								 X"04",X"08",X"80",X"00",
								 X"04",X"08",X"FC",X"00",
								 X"04",X"08",X"C4",X"00",
								 X"04",X"08",X"84",X"00",
								 X"04",X"08",X"86",X"00",
								 X"04",X"18",X"82",X"00",
								 X"02",X"10",X"82",X"00",
								 X"03",X"F0",X"82",X"00",
								 X"00",X"00",X"00",X"00",
								 X"00",X"00",X"00",X"00"),
								----------------------------------------------------
								(X"00",X"00",X"00",X"00", --off
								 X"00",X"01",X"C0",X"60", --15
								 X"00",X"01",X"60",X"F0",
								 X"00",X"01",X"20",X"80",
								 X"00",X"01",X"00",X"80",
								 X"00",X"01",X"00",X"80",
								 X"1F",X"0F",X"E3",X"FC",
								 X"31",X"81",X"00",X"80",
								 X"20",X"81",X"00",X"80",
								 X"20",X"C1",X"00",X"80",
								 X"20",X"41",X"00",X"80",
								 X"10",X"C1",X"00",X"80",
								 X"1F",X"81",X"00",X"80",
								 X"00",X"00",X"00",X"00",
								 X"00",X"00",X"00",X"00",
								 X"00",X"00",X"00",X"00")
								----------------------------------------------------
								);
    ----------------------------------------------------------------------------------------
	type rom16x16 is array (0 to 6, 0 to 31) of std_logic_vector(7 downto 0); 
	constant Font16_1 : rom16x16 :=( -- 16 x 16 / 8 = 32 Bytes (rows x cols = H x W)
								------------------------------------------------------------
								(X"00",X"00",X"00",X"00",X"01",X"80",X"03",X"C0", -- colon (:)
								 X"03",X"C0",X"01",X"80",X"00",X"00",X"00",X"00", -- 0
								 X"00",X"00",X"00",X"00",X"01",X"80",X"03",X"C0",
								 X"03",X"C0",X"01",X"80",X"00",X"00",X"00",X"00"),
								------------------------------------------------------------
								(X"00",X"00",X"00",X"00",X"30",X"00",X"48",X"00", -- deg C
								 X"49",X"F8",X"33",X"FC",X"03",X"0C",X"06",X"00", -- 1
								 X"06",X"00",X"06",X"00",X"06",X"00",X"06",X"00",
								 X"03",X"0C",X"03",X"FC",X"00",X"F8",X"00",X"00"),
								------------------------------------------------------------
								(X"00",X"00",X"30",X"00",X"48",X"00",X"49",X"FC", -- deg F
								 X"31",X"FC",X"01",X"80",X"01",X"80",X"03",X"80", -- 2
								 X"03",X"F8",X"03",X"F8",X"03",X"80",X"03",X"80",
								 X"07",X"00",X"07",X"00",X"07",X"00",X"00",X"00"),
								------------------------------------------------------------
								(X"00",X"00",X"38",X"06",X"44",X"0E",X"44",X"1C", -- percent
								 X"44",X"38",X"38",X"70",X"00",X"E0",X"01",X"C0", -- 3
								 X"03",X"80",X"07",X"00",X"0E",X"1C",X"1C",X"22",
								 X"38",X"22",X"70",X"22",X"60",X"1C",X"00",X"00"),
								------------------------------------------------------------
								(X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- wave(~)
								 X"00",X"00",X"1C",X"00",X"3E",X"00",X"67",X"00", -- 4
								 X"C3",X"86",X"01",X"CC",X"00",X"F8",X"00",X"70",
								 X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								------------------------------------------------------------
								(X"FF",X"FF",X"FF",X"FF",X"7F",X"FE",X"7F",X"FE",
								 X"3F",X"FC",X"3F",X"FC",X"1F",X"F8",X"1F",X"F8",
								 X"0F",X"F0",X"0F",X"F0",X"07",X"E0",X"07",X"E0",
								 X"03",X"C0",X"03",X"C0",X"01",X"80",X"01",X"80"),
								------------------------------------------------------------
								(X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
								 X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
								 X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
								 X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF")
								------------------------------------------------------------
								);
	----------------------------------------------------------------------------------
	-- 111 Contest-1
	type rom128x2 is array(0 to 4,0 to 31) of std_logic_vector(7 downto 0); 
	constant Font128_2 : rom128x2 :=( -- 128 x 2 / 8 = 32 Bytes (rows x cols = H x W)
									 (X"03",X"FF",X"FF",X"FF",X"FC",X"00",X"00",X"00",
									  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
									  X"03",X"FF",X"FF",X"FF",X"FC",X"00",X"00",X"00",
									  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
									 -------------------------------------------------
									 (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",
									  X"FF",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",
									  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",
									  X"FF",X"E0",X"00",X"00",X"00",X"00",X"00",X"00"),
									 -------------------------------------------------
									 (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
									  X"00",X"00",X"00",X"00",X"00",X"7F",X"FF",X"80",
									  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
									  X"00",X"00",X"00",X"00",X"00",X"7F",X"FF",X"80"),
									 -------------------------------------------------
									 (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
									  X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E0",
									  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
									  X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E0"),
									 -------------------------------------------------
									 (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
									  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
									  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
									  X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00")
									 );
    --------------------------------------------------------------------------------
    -- 112 Contest-1 Mode 0 ,2 and 3 (Multi-Characters)
	type rom16x64 is array(0 to 4,0 to 127) of std_logic_vector(7 downto 0); 
	constant Font16_2 : rom16x64 :=( -- 16 x 64 / 8 = 128 Bytes (rows x cols = H x W)
								   -------------------------------------------------
								   -- 0 : Modes:
								   (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",--Modes
									X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
									X"60",X"C0",X"00",X"0C",X"00",X"00",X"0C",X"00",
									X"71",X"C0",X"00",X"0C",X"00",X"00",X"0C",X"00",
									X"7B",X"C0",X"00",X"0C",X"00",X"00",X"00",X"00",
									X"6E",X"C1",X"C0",X"0C",X"7C",X"3F",X"80",X"00",
									X"6E",X"C3",X"E0",X"EC",X"FE",X"7F",X"80",X"00",
									X"64",X"C4",X"11",X"FD",X"C6",X"60",X"00",X"00",
									X"60",X"CC",X"19",X"0D",X"82",X"60",X"00",X"00",
									X"60",X"CC",X"1B",X"0D",X"FE",X"7F",X"00",X"00",
									X"60",X"CC",X"1B",X"0D",X"FC",X"3F",X"80",X"00",
									X"60",X"CC",X"1B",X"0D",X"80",X"01",X"80",X"00",
									X"60",X"C4",X"13",X"0D",X"80",X"01",X"8C",X"00",
									X"60",X"C3",X"E1",X"FC",X"FC",X"7F",X"8C",X"00",
									X"60",X"C1",X"C0",X"FC",X"7E",X"7F",X"00",X"00",
									X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								  --------------------------------------------------
								  -- 1 : Normal
								   (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",--Normal
									X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
									X"60",X"C0",X"00",X"00",X"00",X"00",X"01",X"80",
									X"60",X"C0",X"00",X"00",X"00",X"00",X"01",X"80",
									X"70",X"C3",X"86",X"F6",X"C1",X"83",X"E1",X"80",
									X"78",X"C7",X"C7",X"F7",X"E3",X"E7",X"F1",X"80",
									X"7C",X"CC",X"67",X"87",X"BE",X"E6",X"39",X"80",
									X"6C",X"D8",X"37",X"07",X"1C",X"60",X"19",X"80",
									X"66",X"D8",X"36",X"06",X"18",X"61",X"D9",X"80",
									X"66",X"D8",X"36",X"06",X"18",X"63",X"F9",X"80",
									X"63",X"D8",X"36",X"06",X"18",X"66",X"39",X"80",
									X"63",X"D8",X"36",X"06",X"18",X"66",X"39",X"80",
									X"61",X"CC",X"66",X"06",X"18",X"66",X"39",X"80",
									X"61",X"C7",X"C6",X"06",X"18",X"67",X"F9",X"80",
									X"60",X"C3",X"86",X"06",X"18",X"63",X"F1",X"80",
									X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
                                  --------------------------------------------------
                                  -- 2 : Flash
								  (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", 
								   X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								   X"7F",X"30",X"00",X"00",X"18",X"00",X"00",X"00",
								   X"60",X"30",X"F0",X"1F",X"18",X"00",X"00",X"00",
								   X"60",X"31",X"FC",X"3F",X"98",X"00",X"00",X"00",
								   X"60",X"33",X"0E",X"70",X"18",X"00",X"00",X"00",
								   X"60",X"30",X"06",X"60",X"18",X"00",X"00",X"00",
								   X"7F",X"30",X"F6",X"60",X"1F",X"00",X"00",X"00",
								   X"7F",X"31",X"FE",X"7F",X"1F",X"80",X"00",X"00",
								   X"60",X"33",X"9E",X"3F",X"98",X"C0",X"00",X"00",
								   X"60",X"33",X"0E",X"03",X"98",X"C0",X"00",X"00",
								   X"60",X"33",X"0E",X"01",X"98",X"C0",X"00",X"00",
								   X"60",X"33",X"0E",X"03",X"98",X"C0",X"00",X"00",
								   X"60",X"33",X"FE",X"7F",X"98",X"C0",X"00",X"00",
								   X"60",X"31",X"FC",X"3F",X"18",X"C0",X"00",X"00",
								   X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
								  --------------------------------------------------
								  -- 3 : Speed
								  (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", 
								   X"1F",X"80",X"00",X"00",X"00",X"00",X"60",X"00",
								   X"31",X"C0",X"01",X"F8",X"3F",X"00",X"66",X"00",
								   X"60",X"C7",X"E3",X"FC",X"7F",X"80",X"66",X"00",
								   X"40",X"0F",X"F6",X"06",X"C0",X"C0",X"60",X"00",
								   X"60",X"0C",X"36",X"06",X"C0",X"CF",X"E0",X"00",
								   X"7F",X"0C",X"37",X"FE",X"FF",X"DF",X"E0",X"00",
								   X"3F",X"8C",X"37",X"FC",X"FF",X"98",X"60",X"00",
								   X"01",X"CF",X"F6",X"00",X"C0",X"18",X"60",X"00",
								   X"00",X"CF",X"E6",X"00",X"C0",X"18",X"60",X"00",
								   X"00",X"CC",X"07",X"00",X"C0",X"18",X"60",X"00",
								   X"01",X"CC",X"03",X"FE",X"7F",X"DF",X"E0",X"00",
								   X"3F",X"8C",X"01",X"FC",X"3F",X"8F",X"E6",X"00",
								   X"1F",X"0C",X"00",X"00",X"00",X"00",X"06",X"00",
								   X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
								   X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00"),
								  --------------------------------------------------
								  -- 4 : Moving:
								  (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								   X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
								   X"71",X"C0",X"00",X"00",X"00",X"00",X"06",X"00",
								   X"7B",X"C0",X"00",X"01",X"80",X"00",X"06",X"00",
								   X"6E",X"C0",X"00",X"01",X"80",X"07",X"80",X"00",
								   X"6E",X"C7",X"C0",X"00",X"30",X"0F",X"C0",X"00",
								   X"64",X"CF",X"E6",X"19",X"B7",X"18",X"60",X"00",
								   X"60",X"DC",X"76",X"19",X"BF",X"98",X"60",X"00",
								   X"60",X"D8",X"36",X"19",X"B9",X"D8",X"60",X"00",
								   X"60",X"D8",X"36",X"19",X"B0",X"CF",X"E0",X"00",
								   X"60",X"D8",X"37",X"39",X"B0",X"C7",X"E0",X"00",
								   X"60",X"D8",X"33",X"31",X"B0",X"C0",X"60",X"00",
								   X"60",X"DC",X"73",X"F1",X"B0",X"C0",X"66",X"00",
								   X"60",X"CF",X"E1",X"E1",X"B0",X"CF",X"E6",X"00",
								   X"60",X"C7",X"C0",X"C1",X"B0",X"C7",X"C0",X"00",
								   X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00")
								  );
    --------------------------------------------------------------------------------
    -- 112 Contest-1 Mode 0 ,2 and 3 (Shape Object)
    type rom32x32 is array(0 to 22,0 to 127) of std_logic_vector(7 downto 0); 
	constant Font32_2 : rom32x32 :=( -- 32 x 32 / 8 = 128 Bytes (rows x cols = H x W)
-- 0 : 圓
(
X"00",X"19",X"C8",X"00",X"00",X"AE",X"35",X"00",
X"01",X"E0",X"03",X"80",X"04",X"80",X"00",X"20",
X"0A",X"00",X"00",X"70",X"1C",X"00",X"00",X"28",
X"08",X"00",X"00",X"10",X"20",X"00",X"00",X"04",
X"60",X"00",X"00",X"0E",X"20",X"00",X"00",X"04",
X"40",X"00",X"00",X"06",X"80",X"00",X"00",X"01",
X"40",X"00",X"00",X"03",X"40",X"00",X"00",X"02",
X"80",X"00",X"00",X"02",X"80",X"00",X"00",X"01",
X"80",X"00",X"00",X"01",X"40",X"00",X"00",X"01",
X"40",X"00",X"00",X"02",X"C0",X"00",X"00",X"02",
X"80",X"00",X"00",X"01",X"60",X"00",X"00",X"02",
X"20",X"00",X"00",X"04",X"70",X"00",X"00",X"06",
X"20",X"00",X"00",X"04",X"08",X"00",X"00",X"10",
X"14",X"00",X"00",X"38",X"0E",X"00",X"00",X"50",
X"04",X"00",X"01",X"20",X"01",X"C0",X"07",X"80",
X"00",X"AC",X"75",X"00",X"00",X"13",X"98",X"00"
),
------------------------------------------------
-- 1 : 橢圓
(
X"00",X"09",X"80",X"00",X"00",X"0F",X"F0",X"00",
X"00",X"1F",X"F8",X"00",X"00",X"3F",X"FC",X"00",
X"00",X"7A",X"5F",X"00",X"00",X"70",X"0E",X"00",
X"00",X"78",X"1E",X"00",X"00",X"F0",X"0F",X"00",
X"00",X"F0",X"0F",X"00",X"00",X"F0",X"0F",X"00",
X"00",X"F0",X"0F",X"00",X"00",X"F0",X"0F",X"00",
X"00",X"F0",X"0F",X"00",X"00",X"F0",X"0F",X"00",
X"00",X"F0",X"0F",X"00",X"00",X"F0",X"0F",X"00",
X"00",X"F0",X"0F",X"00",X"00",X"F0",X"0F",X"00",
X"00",X"F0",X"0F",X"00",X"00",X"F0",X"0F",X"00",
X"00",X"F0",X"0F",X"00",X"00",X"F0",X"0F",X"00",
X"00",X"F0",X"0F",X"00",X"00",X"F0",X"0F",X"00",
X"00",X"F0",X"0F",X"00",X"00",X"78",X"1E",X"00",
X"00",X"70",X"0E",X"00",X"00",X"FA",X"5E",X"00",
X"00",X"3F",X"FC",X"00",X"00",X"1F",X"F8",X"00",
X"00",X"0F",X"F0",X"00",X"00",X"01",X"90",X"00"
),
------------------------------------------------
-- 2 : 菱
(
X"00",X"01",X"80",X"00",X"00",X"03",X"C0",X"00",
X"00",X"07",X"A0",X"00",X"00",X"02",X"40",X"00",
X"00",X"04",X"20",X"00",X"00",X"10",X"08",X"00",
X"00",X"28",X"14",X"00",X"00",X"70",X"0E",X"00",
X"00",X"20",X"04",X"00",X"00",X"40",X"02",X"00",
X"01",X"00",X"00",X"80",X"02",X"00",X"00",X"40",
X"07",X"00",X"00",X"E0",X"0A",X"00",X"00",X"50",
X"04",X"00",X"00",X"20",X"08",X"00",X"00",X"00",
X"00",X"00",X"00",X"10",X"04",X"00",X"00",X"20",
X"0A",X"00",X"00",X"50",X"07",X"00",X"00",X"E0",
X"02",X"00",X"00",X"40",X"01",X"00",X"00",X"80",
X"00",X"40",X"02",X"00",X"00",X"20",X"04",X"00",
X"00",X"70",X"0E",X"00",X"00",X"28",X"14",X"00",
X"00",X"10",X"08",X"00",X"00",X"04",X"20",X"00",
X"00",X"02",X"40",X"00",X"00",X"05",X"E0",X"00",
X"00",X"03",X"C0",X"00",X"00",X"01",X"80",X"00"
),
------------------------------------------------
-- 3 : 三角
(
X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
X"00",X"03",X"C0",X"00",X"00",X"01",X"00",X"00",
X"00",X"06",X"20",X"00",X"00",X"02",X"40",X"00",
X"00",X"0C",X"10",X"00",X"00",X"04",X"20",X"00",
X"00",X"18",X"08",X"00",X"00",X"08",X"10",X"00",
X"00",X"30",X"04",X"00",X"00",X"10",X"08",X"00",
X"00",X"60",X"02",X"00",X"00",X"20",X"04",X"00",
X"00",X"80",X"01",X"00",X"00",X"40",X"02",X"00",
X"01",X"00",X"00",X"80",X"00",X"80",X"01",X"00",
X"02",X"00",X"00",X"40",X"01",X"00",X"00",X"80",
X"04",X"00",X"00",X"20",X"02",X"00",X"00",X"40",
X"08",X"00",X"00",X"10",X"04",X"00",X"00",X"20",
X"10",X"00",X"00",X"08",X"08",X"00",X"00",X"10",
X"20",X"00",X"00",X"04",X"10",X"00",X"00",X"08",
X"40",X"00",X"00",X"02",X"20",X"00",X"00",X"04",
X"BF",X"FF",X"FF",X"FD",X"00",X"00",X"00",X"00"
),
------------------------------------------------
-- 4 : 方
(
X"FF",X"FF",X"FF",X"FF",X"80",X"00",X"00",X"01",
X"80",X"00",X"00",X"01",X"80",X"00",X"00",X"01",
X"80",X"00",X"00",X"01",X"80",X"00",X"00",X"01",
X"80",X"00",X"00",X"01",X"80",X"00",X"00",X"01",
X"80",X"00",X"00",X"01",X"80",X"00",X"00",X"01",
X"80",X"00",X"00",X"01",X"80",X"00",X"00",X"01",
X"80",X"00",X"00",X"01",X"80",X"00",X"00",X"01",
X"80",X"00",X"00",X"01",X"80",X"00",X"00",X"01",
X"80",X"00",X"00",X"01",X"80",X"00",X"00",X"01",
X"80",X"00",X"00",X"01",X"80",X"00",X"00",X"01",
X"80",X"00",X"00",X"01",X"80",X"00",X"00",X"01",
X"80",X"00",X"00",X"01",X"80",X"00",X"00",X"01",
X"80",X"00",X"00",X"01",X"80",X"00",X"00",X"01",
X"80",X"00",X"00",X"01",X"80",X"00",X"00",X"01",
X"80",X"00",X"00",X"01",X"80",X"00",X"00",X"01",
X"80",X"00",X"00",X"01",X"FF",X"FF",X"FF",X"FF"
),
------------------------------------------------
-- 5 : 五角
(
X"00",X"01",X"80",X"00",X"00",X"02",X"C0",X"00",
X"00",X"05",X"A0",X"00",X"00",X"12",X"08",X"00",
X"00",X"28",X"1C",X"00",X"00",X"50",X"0A",X"00",
X"01",X"20",X"00",X"80",X"02",X"80",X"01",X"C0",
X"05",X"00",X"00",X"A0",X"12",X"00",X"00",X"08",
X"28",X"00",X"00",X"1C",X"50",X"00",X"00",X"0A",
X"20",X"00",X"00",X"00",X"40",X"00",X"00",X"02",
X"80",X"00",X"00",X"01",X"C0",X"00",X"00",X"02",
X"20",X"00",X"00",X"04",X"40",X"00",X"00",X"02",
X"40",X"00",X"00",X"04",X"10",X"00",X"00",X"08",
X"30",X"00",X"00",X"00",X"20",X"00",X"00",X"0C",
X"08",X"00",X"00",X"18",X"18",X"00",X"00",X"10",
X"10",X"00",X"00",X"08",X"04",X"00",X"00",X"10",
X"04",X"00",X"00",X"20",X"08",X"00",X"00",X"10",
X"06",X"00",X"00",X"20",X"02",X"00",X"00",X"40",
X"04",X"00",X"00",X"20",X"07",X"FF",X"FF",X"C0"
),
------------------------------------------------
-- 6 : 六角
(
X"00",X"00",X"00",X"00",X"01",X"7F",X"FF",X"40",
X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",
X"02",X"00",X"00",X"00",X"02",X"00",X"00",X"70",
X"0C",X"00",X"00",X"10",X"04",X"00",X"00",X"20",
X"18",X"00",X"00",X"08",X"08",X"00",X"00",X"10",
X"30",X"00",X"00",X"04",X"10",X"00",X"00",X"08",
X"60",X"00",X"00",X"02",X"20",X"00",X"00",X"04",
X"80",X"00",X"00",X"01",X"40",X"00",X"00",X"02",
X"40",X"00",X"00",X"02",X"80",X"00",X"00",X"01",
X"20",X"00",X"00",X"04",X"40",X"00",X"00",X"02",
X"10",X"00",X"00",X"08",X"20",X"00",X"00",X"04",
X"08",X"00",X"00",X"18",X"10",X"00",X"00",X"08",
X"04",X"00",X"00",X"30",X"0E",X"00",X"00",X"10",
X"00",X"00",X"00",X"20",X"07",X"00",X"00",X"00",
X"00",X"00",X"00",X"40",X"03",X"80",X"00",X"80",
X"00",X"7F",X"FF",X"C0",X"00",X"00",X"00",X"00"
),
------------------------------------------------
-- 7 : 倒三角
(
X"00",X"00",X"00",X"00",X"BF",X"FF",X"FF",X"FD",
X"20",X"00",X"00",X"04",X"40",X"00",X"00",X"02",
X"10",X"00",X"00",X"08",X"20",X"00",X"00",X"04",
X"08",X"00",X"00",X"10",X"10",X"00",X"00",X"08",
X"04",X"00",X"00",X"20",X"08",X"00",X"00",X"10",
X"02",X"00",X"00",X"40",X"04",X"00",X"00",X"20",
X"01",X"00",X"00",X"80",X"02",X"00",X"00",X"40",
X"00",X"80",X"01",X"00",X"01",X"00",X"00",X"80",
X"00",X"40",X"02",X"00",X"00",X"80",X"01",X"00",
X"00",X"20",X"04",X"00",X"00",X"40",X"06",X"00",
X"00",X"10",X"08",X"00",X"00",X"20",X"0C",X"00",
X"00",X"08",X"10",X"00",X"00",X"10",X"18",X"00",
X"00",X"04",X"20",X"00",X"00",X"08",X"30",X"00",
X"00",X"02",X"40",X"00",X"00",X"04",X"60",X"00",
X"00",X"00",X"80",X"00",X"00",X"03",X"C0",X"00",
X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00"
),
------------------------------------------------
-- 8 : 八角
(
X"00",X"7F",X"FE",X"00",X"00",X"80",X"01",X"00",
X"01",X"00",X"00",X"80",X"02",X"00",X"00",X"40",
X"04",X"00",X"00",X"20",X"08",X"00",X"00",X"10",
X"10",X"00",X"00",X"08",X"20",X"00",X"00",X"04",
X"40",X"00",X"00",X"02",X"80",X"00",X"00",X"01",
X"80",X"00",X"00",X"01",X"80",X"00",X"00",X"01",
X"80",X"00",X"00",X"01",X"80",X"00",X"00",X"01",
X"80",X"00",X"00",X"01",X"80",X"00",X"00",X"01",
X"80",X"00",X"00",X"01",X"80",X"00",X"00",X"01",
X"80",X"00",X"00",X"01",X"80",X"00",X"00",X"01",
X"80",X"00",X"00",X"01",X"80",X"00",X"00",X"01",
X"80",X"00",X"00",X"01",X"80",X"00",X"00",X"02",
X"40",X"00",X"00",X"04",X"20",X"00",X"00",X"08",
X"10",X"00",X"00",X"10",X"08",X"00",X"00",X"20",
X"04",X"00",X"00",X"40",X"02",X"00",X"00",X"80",
X"01",X"00",X"01",X"00",X"00",X"FF",X"FE",X"00"
),
------------------------------------------------
-- 9 : 長方形
(
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"FF",X"FF",X"FF",X"FF",X"80",X"00",X"00",X"01",
X"80",X"00",X"00",X"01",X"80",X"00",X"00",X"01",
X"80",X"00",X"00",X"01",X"80",X"00",X"00",X"01",
X"80",X"00",X"00",X"01",X"80",X"00",X"00",X"01",
X"80",X"00",X"00",X"01",X"80",X"00",X"00",X"01",
X"80",X"00",X"00",X"01",X"FF",X"FF",X"FF",X"FF",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"
),
------------------------------------------------
-- 10 : 滿圓
(
X"00",X"1B",X"C8",X"00",X"00",X"BF",X"FD",X"00",
X"01",X"FF",X"FF",X"80",X"07",X"FF",X"FF",X"A0",
X"0F",X"FF",X"FF",X"F0",X"1F",X"FF",X"FF",X"F8",
X"0F",X"FF",X"FF",X"F8",X"3F",X"FF",X"FF",X"FC",
X"7F",X"FF",X"FF",X"FE",X"3F",X"FF",X"FF",X"FC",
X"7F",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",
X"7F",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FE",
X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
X"7F",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FE",
X"FF",X"FF",X"FF",X"FF",X"7F",X"FF",X"FF",X"FE",
X"3F",X"FF",X"FF",X"FC",X"7F",X"FF",X"FF",X"FE",
X"3F",X"FF",X"FF",X"FC",X"1F",X"FF",X"FF",X"F0",
X"1F",X"FF",X"FF",X"F8",X"0F",X"FF",X"FF",X"F0",
X"05",X"FF",X"FF",X"E0",X"01",X"FF",X"FF",X"80",
X"00",X"BF",X"FD",X"00",X"00",X"13",X"D8",X"00"
),
------------------------------------------------
-- 11 : 滿橢圓
(
X"00",X"0B",X"D0",X"00",X"00",X"0F",X"F0",X"00",
X"00",X"1F",X"F8",X"00",X"00",X"3F",X"FC",X"00",
X"00",X"FF",X"FF",X"00",X"00",X"7F",X"FE",X"00",
X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",
X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",
X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",
X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",
X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",
X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",
X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",
X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",
X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",
X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",
X"00",X"7F",X"FE",X"00",X"00",X"FF",X"FF",X"00",
X"00",X"3F",X"FC",X"00",X"00",X"1F",X"F8",X"00",
X"00",X"0F",X"F0",X"00",X"00",X"0B",X"D0",X"00"
),
------------------------------------------------
-- 12 : 滿菱
(
X"00",X"01",X"80",X"00",X"00",X"03",X"C0",X"00",
X"00",X"07",X"E0",X"00",X"00",X"03",X"E0",X"00",
X"00",X"07",X"E0",X"00",X"00",X"1F",X"F8",X"00",
X"00",X"3F",X"FC",X"00",X"00",X"7F",X"FE",X"00",
X"00",X"7F",X"FE",X"00",X"00",X"7F",X"FE",X"00",
X"01",X"FF",X"FF",X"80",X"03",X"FF",X"FF",X"C0",
X"07",X"FF",X"FF",X"E0",X"0F",X"FF",X"FF",X"F0",
X"07",X"FF",X"FF",X"E0",X"0F",X"FF",X"FF",X"F0",
X"0F",X"FF",X"FF",X"F0",X"07",X"FF",X"FF",X"E0",
X"0F",X"FF",X"FF",X"F0",X"07",X"FF",X"FF",X"E0",
X"03",X"FF",X"FF",X"C0",X"01",X"FF",X"FF",X"80",
X"00",X"7F",X"FE",X"00",X"00",X"7F",X"FE",X"00",
X"00",X"7F",X"FE",X"00",X"00",X"3F",X"FC",X"00",
X"00",X"1F",X"F8",X"00",X"00",X"07",X"E0",X"00",
X"00",X"07",X"C0",X"00",X"00",X"07",X"E0",X"00",
X"00",X"03",X"C0",X"00",X"00",X"01",X"80",X"00"
),
------------------------------------------------
-- 13 : 滿三角
(
X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
X"00",X"01",X"40",X"00",X"00",X"00",X"80",X"00",
X"00",X"02",X"A0",X"00",X"00",X"01",X"C0",X"00",
X"00",X"07",X"D0",X"00",X"00",X"07",X"F0",X"00",
X"00",X"0F",X"E8",X"00",X"00",X"0F",X"F8",X"00",
X"00",X"1F",X"F4",X"00",X"00",X"1F",X"FE",X"00",
X"00",X"1F",X"FC",X"00",X"00",X"7F",X"FF",X"00",
X"00",X"3F",X"FE",X"00",X"00",X"FF",X"FE",X"80",
X"00",X"7F",X"FF",X"00",X"01",X"FF",X"FF",X"40",
X"00",X"FF",X"FF",X"C0",X"03",X"FF",X"FF",X"A0",
X"03",X"FF",X"FF",X"E0",X"05",X"FF",X"FF",X"D0",
X"07",X"FF",X"FF",X"F8",X"0F",X"FF",X"FF",X"E0",
X"1F",X"FF",X"FF",X"FC",X"0F",X"FF",X"FF",X"F8",
X"3F",X"FF",X"FF",X"FA",X"1F",X"FF",X"FF",X"FC",
X"5F",X"FF",X"FF",X"FD",X"3F",X"FF",X"FF",X"FE",
X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00"
),
------------------------------------------------
-- 14 : 滿方
(
X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF"
),
------------------------------------------------
-- 15 : 滿五角
(
X"00",X"01",X"00",X"00",X"00",X"03",X"C0",X"00",
X"00",X"0F",X"F0",X"00",X"00",X"13",X"E8",X"00",
X"00",X"77",X"F6",X"00",X"00",X"FF",X"FF",X"00",
X"01",X"3F",X"FC",X"80",X"06",X"7F",X"FE",X"60",
X"0F",X"FF",X"FF",X"F0",X"1B",X"FF",X"FF",X"F8",
X"27",X"FF",X"FF",X"E6",X"FF",X"FF",X"FF",X"FF",
X"FF",X"FF",X"FF",X"FE",X"7F",X"FF",X"FF",X"FE",
X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
X"3F",X"FF",X"FF",X"FC",X"5F",X"FF",X"FF",X"FE",
X"5F",X"FF",X"FF",X"FE",X"1F",X"FF",X"FF",X"F8",
X"2F",X"FF",X"FF",X"FC",X"3F",X"FF",X"FF",X"FC",
X"1F",X"FF",X"FF",X"F0",X"1F",X"FF",X"FF",X"F8",
X"17",X"FF",X"FF",X"F8",X"0F",X"FF",X"FF",X"F8",
X"07",X"FF",X"FF",X"E0",X"0B",X"FF",X"FF",X"F0",
X"07",X"FF",X"FF",X"D0",X"03",X"FF",X"FF",X"C0",
X"05",X"FF",X"FF",X"E0",X"07",X"FF",X"FF",X"C0"
),
------------------------------------------------
-- 16 : 滿六角
(
X"00",X"00",X"00",X"00",X"01",X"FF",X"FF",X"C0",
X"01",X"FF",X"FF",X"00",X"03",X"FF",X"FF",X"C0",
X"07",X"FF",X"FF",X"A0",X"07",X"FF",X"FF",X"F0",
X"0F",X"FF",X"FF",X"D0",X"0F",X"FF",X"FF",X"F8",
X"1F",X"FF",X"FF",X"E8",X"1F",X"FF",X"FF",X"F8",
X"3F",X"FF",X"FF",X"F4",X"1F",X"FF",X"FF",X"FA",
X"7F",X"FF",X"FF",X"FA",X"3F",X"FF",X"FF",X"FD",
X"FF",X"FF",X"FF",X"FD",X"7F",X"FF",X"FF",X"FC",
X"3F",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",
X"5F",X"FF",X"FF",X"FC",X"7F",X"FF",X"FF",X"FE",
X"2F",X"FF",X"FF",X"FA",X"3F",X"FF",X"FF",X"F4",
X"17",X"FF",X"FF",X"F4",X"1F",X"FF",X"FF",X"F8",
X"0B",X"FF",X"FF",X"E8",X"0F",X"FF",X"FF",X"F0",
X"05",X"FF",X"FF",X"D0",X"07",X"FF",X"FF",X"E0",
X"02",X"FF",X"FF",X"E0",X"01",X"FF",X"FF",X"C0",
X"01",X"7F",X"FF",X"80",X"00",X"00",X"00",X"00"
),
------------------------------------------------
-- 17 : 滿倒三角
(
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"70",X"FF",X"80",X"00",X"BF",X"FF",X"FF",X"FF",
X"7F",X"FF",X"FF",X"FD",X"5F",X"FF",X"FF",X"FA",
X"2F",X"FF",X"FF",X"FC",X"07",X"FF",X"FF",X"F4",
X"1F",X"FF",X"FF",X"E8",X"0F",X"FF",X"FF",X"E8",
X"0B",X"FF",X"FF",X"D0",X"07",X"FF",X"FF",X"80",
X"04",X"FF",X"FF",X"A0",X"03",X"FF",X"FF",X"40",
X"00",X"FF",X"FF",X"00",X"01",X"FF",X"FE",X"80",
X"00",X"BF",X"FC",X"00",X"00",X"FF",X"FF",X"00",
X"00",X"1F",X"FA",X"00",X"00",X"5F",X"FC",X"00",
X"00",X"3F",X"FC",X"00",X"00",X"0F",X"E0",X"00",
X"00",X"17",X"F8",X"00",X"00",X"07",X"D0",X"00",
X"00",X"0B",X"F0",X"00",X"00",X"03",X"A0",X"00",
X"00",X"05",X"80",X"00",X"00",X"03",X"C0",X"00",
X"00",X"02",X"00",X"00",X"00",X"01",X"80",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"
),
------------------------------------------------
-- 18 : 滿八角
(
X"00",X"7F",X"FE",X"00",X"00",X"FF",X"FF",X"00",
X"01",X"FF",X"FF",X"80",X"03",X"FF",X"FF",X"C0",
X"07",X"FF",X"FF",X"E0",X"0F",X"FF",X"FF",X"F0",
X"1F",X"FF",X"FF",X"F8",X"3F",X"FF",X"FF",X"FC",
X"7F",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",
X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",
X"7F",X"FF",X"FF",X"FC",X"3F",X"FF",X"FF",X"F8",
X"1F",X"FF",X"FF",X"F0",X"0F",X"FF",X"FF",X"E0",
X"07",X"FF",X"FF",X"C0",X"03",X"FF",X"FF",X"80",
X"01",X"FF",X"FF",X"00",X"00",X"FF",X"FE",X"00"
),
------------------------------------------------
-- 19 : 滿長方
(
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"
),
------------------------------------------------
-- 20 : 空白
(
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"
),
------------------------------------------------
-- 21 : WIFI
(
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"0F",X"F8",X"00",X"00",X"3F",X"FC",X"00",
X"01",X"FF",X"FF",X"80",X"03",X"FF",X"FF",X"E0",
X"0F",X"F0",X"0B",X"F0",X"0F",X"80",X"01",X"F0",
X"3C",X"00",X"00",X"78",X"3C",X"1F",X"F8",X"3C",
X"70",X"7F",X"FE",X"1E",X"70",X"7F",X"FE",X"0E",
X"71",X"FF",X"7F",X"8C",X"03",X"F0",X"0F",X"80",
X"07",X"E0",X"07",X"E0",X"07",X"80",X"01",X"E0",
X"07",X"0F",X"F0",X"E0",X"06",X"1F",X"F8",X"60",
X"00",X"3F",X"FC",X"00",X"00",X"7F",X"FE",X"00",
X"00",X"74",X"3E",X"00",X"00",X"70",X"06",X"00",
X"00",X"60",X"02",X"00",X"00",X"00",X"00",X"00",
X"00",X"03",X"C0",X"00",X"00",X"07",X"E0",X"00",
X"00",X"07",X"E0",X"00",X"00",X"07",X"E0",X"00",
X"00",X"07",X"E0",X"00",X"00",X"03",X"C0",X"00",
X"00",X"03",X"C0",X"00",X"00",X"00",X"00",X"00"
),
------------------------------------------------
-- 22 : 滿直長方
(
X"00",X"3F",X"FC",X"00",X"00",X"3F",X"FC",X"00",
X"00",X"3F",X"FC",X"00",X"00",X"3F",X"FC",X"00",
X"00",X"3F",X"FC",X"00",X"00",X"3F",X"FC",X"00",
X"00",X"3F",X"FC",X"00",X"00",X"3F",X"FC",X"00",
X"00",X"3F",X"FC",X"00",X"00",X"3F",X"FC",X"00",
X"00",X"3F",X"FC",X"00",X"00",X"3F",X"FC",X"00",
X"00",X"3F",X"FC",X"00",X"00",X"3F",X"FC",X"00",
X"00",X"3F",X"FC",X"00",X"00",X"3F",X"FC",X"00",
X"00",X"3F",X"FC",X"00",X"00",X"3F",X"FC",X"00",
X"00",X"3F",X"FC",X"00",X"00",X"3F",X"FC",X"00",
X"00",X"3F",X"FC",X"00",X"00",X"3F",X"FC",X"00",
X"00",X"3F",X"FC",X"00",X"00",X"3F",X"FC",X"00",
X"00",X"3F",X"FC",X"00",X"00",X"3F",X"FC",X"00",
X"00",X"3F",X"FC",X"00",X"00",X"3F",X"FC",X"00",
X"00",X"3F",X"FC",X"00",X"00",X"3F",X"FC",X"00",
X"00",X"3F",X"FC",X"00",X"00",X"3F",X"FC",X"00"
));
--**********************************************************************************
begin
-- System Connections
	BL_tft <= '1'; -- Back-Light On
--	BL_tft <= '0'; -- Back-Light Off
--**********************************************************************************
x1 : block
    -- RGB TFT LCD SPI FSM's Signals
	type   states is ( s0, s1, s2, s3, s4, s5, s6, s7, s8, s9,s10,s11,s12,s13,s14,
					  s15,s16,s17,s18,s19,s20,s21,s22,s23,s24,s25,s26,s27,s28,s29,
					  s30,s31,s32,s33,s34,s35,s36);
	signal ps,ns  : states;
	--------------------------------------------------------------------------------
	-- ST7735 指令 & 資料表格式 :
	type ROM is array (0 to 84) of std_logic_vector(7 Downto 0);
	-- ST7735 初始化指令表 :
	constant cmd_ROM:ROM :=(--------------------------------------------------------
							X"11", -- 00 SLPOUT    : Sleep out & Booster on 
							--------------------------------------------------------
                            X"B1", -- 01 FRMCTR1   : Frame Rate Control-1
							X"05", -- 02 Payload 1
							X"3C", -- 03 Payload 2
							X"3C", -- 04 Payload 3
							--------------------------------------------------------
							X"B2", -- 05 FRMCTR2   : Frame Rate Control-2
							X"05", -- 06 Payload 1
							X"3C", -- 07 Payload 2
							X"3C", -- 08 Payload 3
							--------------------------------------------------------
							X"B3", -- 09 FRMCTR3   : Frame Rate Control-3
							X"05", -- 10 Payload 1
							X"3C", -- 11 Payload 2
							X"3C", -- 12 Payload 3
							X"05", -- 13 Payload 4
							X"3C", -- 14 Payload 5
							X"3C", -- 15 Payload 6
							--------------------------------------------------------
						    X"B4", -- 16 INVCTR   : Display Inversion Control
						    X"03", -- 17 Payload 1
						    --------------------------------------------------------
                            X"C0", -- 18 PWCTR1   : Power Control-1
							X"28", -- 19 Payload 1
							X"08", -- 20 Payload 2
--							X"04", --    Payload 3 /!\
							--------------------------------------------------------
							X"C1", -- 21 PWCTR2   : Power Control-2
							X"C0", -- 22 Payload 1
							--------------------------------------------------------
							X"C2", -- 23 PWCTR3   : Power Control-3
							X"0D", -- 24 Payload 1
							X"00", -- 25 Payload 2
							--------------------------------------------------------
							X"C3", -- 26 PWCTR4   : Power Control-4
							X"8D", -- 27 Payload 1
							X"2A", -- 28 Payload 2
							--------------------------------------------------------
							X"C4", -- 29 PWCTR5   : Power Control-5
							X"8D", -- 30 Payload 1
							X"EE", -- 31 Payload 2
							--------------------------------------------------------
							X"C5", -- 32 VMCTR1   : VCOM Control-1 
							X"18", -- 33 Payload 1 or X"18"
							X"1A", -- 34 Payload 2 /!\
							--------------------------------------------------------
							X"36", -- 35 MADCTL    : Memory data access control
							X"C0", -- 36 Payload 1 : MY-MX-MV-ML-RGB-MH-x-x
								   --                1  1  0  0   0  0  0 0
								   --    Mirror-Y ,  Mirror-X
							--------------------------------------------------------
							X"E0", -- 37 GAMCTRP1 : Gamma adjustment + polarity
							X"04", -- 38 Payload  1
							X"22", -- 39 Payload  2
							X"07", -- 40 Payload  3
							X"0A", -- 41 Payload  4
							X"2E", -- 42 Payload  5
							X"30", -- 43 Payload  6
							X"25", -- 44 Payload  7
							X"2A", -- 45 Payload  8
							X"28", -- 46 Payload  9
							X"26", -- 47 Payload 10
							X"2E", -- 48 Payload 11
							X"3A", -- 49 Payload 12
							X"00", -- 50 Payload 13
							X"01", -- 51 Payload 14
							X"03", -- 52 Payload 15
							X"13", -- 53 Payload 16
                            --------------------------------------------------------
							X"E1", -- 54 GAMCTRN1 : Gamma adjustment - polarity
							X"04", -- 55 Payload  1
							X"16", -- 56 Payload  2
							X"06", -- 57 Payload  3
							X"0D", -- 58 Payload  4
							X"2D", -- 59 Payload  5
							X"26", -- 60 Payload  6
							X"23", -- 61 Payload  7
							X"27", -- 62 Payload  8
							X"27", -- 63 Payload  9
							X"25", -- 64 Payload 10
							X"2D", -- 65 Payload 11
							X"3B", -- 66 Payload 12
							X"00", -- 67 Payload 13
							X"01", -- 68 Payload 14
							X"04", -- 69 Payload 15
							X"13", -- 70 Payload 16
						    --------------------------------------------------------
							X"3A", -- 71 COLMOD    : Interface Pixel Format
							X"05", -- 72 Payload 1 : 16 Bits / Pixel
							--------------------------------------------------------
							X"29", -- 73 DISPON    : Display On 
							--------------------------------------------------------
							X"2A", -- 74 CASET     : Column Address Set
							X"00", -- 75 Payload 1 ; XS = 0x0002 =   2
							X"02", -- 76 Payload 2
							X"00", -- 77 Payload 3 ; XE = 0x0081 = 129
							X"81", -- 78 Payload 4
							--------------------------------------------------------
							X"2B", -- 79 RASET     : Row    Address Set
							X"00", -- 80 Payload 1 ; YS = 0x0001 =   1
							X"01", -- 81 Payload 2
							X"00", -- 82 Payload 3 ; YE = 0x00A0 = 160
							X"A0", -- 83 Payload 4
							--------------------------------------------------------
							X"2C"  -- 84 RAMWR    : RAM Write (....) CS = 0
							--------------------------------------------------------
						   );
    --------------------------------------------------------------------------------
	type table is array (0 to 84) of std_logic;
	constant DC_table:table :=(	----------------------------------------------------
							'0', -- 00  SLPOUT  : Sleep out & Booster on
							--------------------------------------------------------
                            '0', -- 01  FRMCTR1 : Frame Rate Control-1
							'1', -- 02
							'1', -- 03
							'1', -- 04
							--------------------------------------------------------
							'0', -- 05  FRMCTR2 : Frame Rate Control-2
							'1', -- 06
							'1', -- 07
							'1', -- 08
							--------------------------------------------------------
							'0', -- 09  FRMCTR3 : Frame Rate Control-3
							'1', -- 10
							'1', -- 11
							'1', -- 12
							'1', -- 13
							'1', -- 14
							'1', -- 15
							--------------------------------------------------------
							'0', -- 16  INVCTR : Display Inversion Control
							'1', -- 17
						    --------------------------------------------------------
							'0', -- 18
							'1', -- 19
							'1', -- 20
--							'1', --     /!\
							--------------------------------------------------------
							'0', -- 21
							'1', -- 22
							--------------------------------------------------------
							'0', -- 23
							'1', -- 24
							'1', -- 25
							--------------------------------------------------------
							'0', -- 26
							'1', -- 27
							'1', -- 28
							--------------------------------------------------------
							'0', -- 29
							'1', -- 30
							'1', -- 31
							--------------------------------------------------------
							'0', -- 32  VMCTR1 : VCOM Control-1 
							'1', -- 33
							'1', -- 34  /!\
							--------------------------------------------------------
							'0', -- 35  MADCTL : Memory data access control
							'1', -- 36           MY-MX-MV-ML-RGB-MH-x-x
							--------------------------------------------------------
							'0', -- 37  GAMCTRP1 : Gamma adjustment + polarity
							'1', -- 38
							'1', -- 39
							'1', -- 40
							'1', -- 41
							'1', -- 42
							'1', -- 43
							'1', -- 44
							'1', -- 45
							'1', -- 46
							'1', -- 47
							'1', -- 48
							'1', -- 49
							'1', -- 50
							'1', -- 51
							'1', -- 52
							'1', -- 53
							--------------------------------------------------------
							'0', -- 54  GAMCTRN1 : Gamma adjustment - polarity
							'1', -- 55
							'1', -- 56
							'1', -- 57
							'1', -- 58
							'1', -- 59
							'1', -- 60
							'1', -- 61
							'1', -- 62
							'1', -- 63
							'1', -- 64
							'1', -- 65
							'1', -- 66
							'1', -- 67
							'1', -- 68
							'1', -- 69
							'1', -- 70
						    -------------------------------------------------------- 
							'0', -- 71  COLMOD : Interface Pixel Format
							'1', -- 72
							--------------------------------------------------------
							'0', -- 73 DISPON
							--------------------------------------------------------
							'0', -- 74  CASET : Column Address Set
							'1', -- 75
							'1', -- 76
							'1', -- 77
							'1', -- 78
							--------------------------------------------------------
							'0', -- 79  RASET : Row Address Set
							'1', -- 80
							'1', -- 81
							'1', -- 82
							'1', -- 83
							--------------------------------------------------------
							'0'  -- 84  RAMWR : RAM Write (....) CS = 0
							--------------------------------------------------------
							);
	--------------------------------------------------------------------------------
	type RAM1 is array (0 to 10) of std_logic_vector(7 Downto 0);
	constant cmd_RAM : RAM1 :=( ----------------------------------------------------
								X"2A", -- 00 CASET     : Column Address Set
								X"00", -- 01 Payload 1 ; X1 = 0x0002 =   2
								X"02", -- 02 Payload 2
								X"00", -- 03 Payload 3 ; X2 = 0x0081 = 129
								X"81", -- 04 Payload 4
								----------------------------------------------------
								X"2B", -- 05 RASET     : Row    Address Set
								X"00", -- 06 Payload 1 ; Y1 = 0x0001 =   1
								X"01", -- 07 Payload 2
								X"00", -- 08 Payload 3 ; Y2 = 0x00A0 = 160
								X"A0", -- 09 Payload 4
								----------------------------------------------------
								X"2C"  -- 10 RAMWR     : RAM Write (....) cs = 0
								----------------------------------------------------
							  );
	signal cmd_RAM1 : RAM1;
    --------------------------------------------------------------------------------
	type RAM2 is array (0 to 10) of std_logic;
	constant DC_RAM : RAM2 :=(------------------------------------------------------
							  '0', -- 00 CASET : Column Address Set
							  '1', -- 01
							  '1', -- 02
							  '1', -- 03
							  '1', -- 04
							  ------------------------------------------------------
							  '0', -- 05 RASET : Row    Address Set
							  '1', -- 06
							  '1', -- 07
							  '1', -- 08
							  '1', -- 09
							  ------------------------------------------------------
							  '0'  -- 10 RAMWR : RAM Write (....) cs = 0
							 -------------------------------------------------------
                             );
	signal DC_RAM1 : RAM2;
------------------------------------------------------------------------------------
begin
	--------------------------------------------------------------------------------
	-- Two Processes FSM
	--------------------------------------------------------------------------------
	-- (1) State changing
	process(clk,rst) -- Sensitivity List 
	begin
		if(rst = '0')then -- Initializations (Asynchronous Reset)
			ps <= s0;
		elsif(clk'event and clk = '1')then -- Positive-Edge Trigger (20nS)
			ps <= ns;
		end if;
	end process;
	--------------------------------------------------------------------------------
	-- (2) Individual state excution sequence
	process(clk,rst) -- Sensitivity List
		variable cnt   : integer ;                   -- 32 bits
		variable cnt0  : integer range 0 to     160; --  8 bits
		variable cnt1  : integer range 0 to     128; --  8 bits
		variable cnt2  : integer range 0 to      15; --  4 bits
		variable cnt3  : integer range 0 to      31; --  5 bits
		variable index : integer range 0 to   20480; -- 15 bits
		variable cnt_r : integer range 0 to     128; --  8 bits
	--------------------------------------------------------------------------------
	begin
		if(rst = '0')then      -- Initializations (Asynchronous Reset)
			rst_tft    <= '1'; -- Reset Disable
			cs         <= '1'; -- CS    Disable
			dc		   <= '0'; -- Command
			scl 	   <= '0'; -- Idled State
			sda 	   <= '0';
			ns  	   <= s0;
			bf_out     <= '1';  -- 1 : Busy
			flag_init  <= "01"; -- Entry RGB TFT LCD Initializations
			flag_start <= '0';
			for i in 0 to 10 loop
				cmd_RAM1(i) <= cmd_RAM(i);
				DC_RAM1(i)  <= DC_RAM(i);
			end loop;
        elsif(clk'event and clk = '0')then -- Negative-Edge Trigger (20nS)
			------------------------------------------------------------------------
			-- 1. RGB TFT LCD Initialization Settings
			------------------------------------------------------------------------
			if(flag_init = "01")then -- 20nS
				flag_init  <= "10";
				flag_start <= '0';
				bf_out     <= '1'; -- 1 : busy
				index      := 0;
				cnt        := 0;
				ns         <= s0; 
			------------------------------------------------------------------------
			-- 2. RGB TFT LCD Initialization Sequences
			------------------------------------------------------------------------
			elsif(flag_init = "10" and tft_lcd_p = '1')then -- 100nS
				case ps is -- 100nS
					----------------------------------------------------------------
					-- (1) ST7735 Reset Sequences
					----------------------------------------------------------------
					when s0 => -- rst_tft holds High for 1mS
						rst_tft <= '1'; -- Reset Disable
						cs      <= '1'; -- CS    Disable
						dc      <= '0'; -- Command
						scl     <= '0'; -- Idled State
						sda     <= '0';
						if(cnt < 1E4)then
							cnt := cnt + 1;
							ns  <= s0;
						else
							cnt := 0;
							ns  <= s1;
						end if;
					when s1 =>	-- rst_tft holds Low for 1mS
						rst_tft <= '0'; -- Reset ST7735
						cs      <= '1'; -- CS    Disable
						dc      <= '0'; -- Command
						scl     <= '0'; -- Idled State
						sda     <= '0';
						if(cnt < 1E4)then
							cnt := cnt + 1;
							ns  <= s1;
						else
							cnt := 0;
							ns  <= s2;
						end if;
					when s2 => -- rst_tft holds High for 120mS
						rst_tft <= '1'; -- Reset Disable
						cs      <= '1'; -- CS    Disable
						dc      <= '0'; -- Command
						scl     <= '0'; -- Idled State
						sda     <= '0';
						if(cnt < 12E5)then -- 100nS * 1200000 = 120mS 
							cnt := cnt + 1;
							ns  <= s2;
						else
							cnt := 0;
							ns  <= s3;
						end if;
					----------------------------------------------------------------
					-- (2) Sleep out & Booster on
					----------------------------------------------------------------
					when s3 =>  
						code    <= cmd_ROM(0); -- 0x"11"
						rst_tft <= '1'; -- Reset Disable
						cs      <= '1'; -- CS    Disable
						dc      <= '0'; -- Command 
						scl     <= '0'; -- Idled State
						sda     <= '0';
						cnt     := 8;   -- 8 Bits                    
						ns      <= s4;
					when s4 =>
						cs  <= '0'; -- CS Falling-Edge Trigger : Start Sequence
						scl <= '0';
						if(code(cnt - 1) = '0')then -- MSB First Tx
							sda <= '0';
						else
							sda <= '1';
						end if;
						ns <= s5;
					when s5 => 
						scl <= '1'; -- Positive-Edge Trigger
						if(cnt > 1)then 
							cnt := cnt - 1;
							ns  <= s4;
						else
							cnt := 0;
							ns  <= s6;
						end if;
					when s6 =>
						scl <= '0'; -- Idled State
						sda <= '0';
						ns  <= s7;
					when s7 =>
						cs  <= '1'; -- Rising-Edge Trigger : Stop Sequence
						dc  <= '0'; -- Command                         
						ns  <= s8;                   
					when s8 => -- Waiting 120 mS
						if(cnt < 12E5)then
							cnt := cnt + 1;
							ns  <= s8;
						else
							cnt := 0;
							ns  <= s9;
						end if;
					----------------------------------------------------------------
					-- (3) Two-Loops : Initial Command and Parameters
					----------------------------------------------------------------
					when s9 => -- Outer Loop Parameters Setting
						index :=  1;
						cs    <= '1'; -- CS Disable
						scl   <= '0';
						sda   <= '0'; 
						ns    <= s10;
					when s10 => -- Outer Loop (Inner Loop Parameters Setting)
						code <= cmd_ROM(index);
						dc   <= DC_table(index); -- Command or Parameter 
						cnt2 := 8;               -- 8 Bits              
						ns   <= s11;
					when s11 => -- Inner Loop (Parameters Setting)
						cs   <= '0'; -- CS Falling-Edge Trigger : Start Sequence
						scl  <= '0';
						if(code(cnt2 - 1) = '0')then -- MSB First Tx
							sda <= '0';
						else
							sda <= '1';
						end if;
						ns <= s12;                   
					when s12 =>
						scl <= '1'; -- Positive-Edge Trigger
						if(cnt2 > 1)then 
							cnt2 := cnt2 - 1;
							ns   <= s11; -- Return to Inner Loop
						else 
							ns  <= s13;
						end if; 
					when s13 =>
						scl <= '0';
						sda <= '0';
						if(index < 84)then -- 84 : RAMWR (....) , CS = 0
							index := index + 1;
							ns    <= s10; -- Return to Outer Loop
						else
							cnt2 := 8;   -- 8 Bits
							ns   <= s14; -- /!\ 
						end if;
					----------------------------------------------------------------
					-- (4) Setting 128 x 160 Pixels Color
					----------------------------------------------------------------
					when s14 =>
						dc     <= '1'; -- Data
						scl    <= '0';
						sda    <= '0';
						color  <= X"FFFF"; -- RGB : 5-6-5 -> 16 Bits (White)
						index  := 0;       -- RGB Color Start index
						cnt3   := 16;      -- 16 Bits (R-G-B : 5-6-5)
						ns     <= s15;
					----------------------------------------------------------------
					when s15 => -- Outer Loop
						scl   <= '0';
						sda   <= '0';
						ns    <= s16;      
					when s16 => -- Inner Loop 
						scl  <= '0';
						if(color(cnt3 - 1) = '0')then -- MSB First Tx
							sda <= '0';
						else
							sda <= '1';
						end if;
						ns <= s17;
					when s17 =>
						scl <= '1'; -- Positive-Edge Trigger
						if(cnt3 > 1)then 
							cnt3 := cnt3 - 1;
							ns   <= s16; -- Inner Loop
						else 
							ns <= s18;
						end if;                   
					when s18 =>
						scl <= '0';
						sda <= '0';
						if(index < 20480)then -- 160 x 128 = 20480 Pixels
							index := index + 1;
							cnt3  := 16;
							color <= X"0000"; -- Black
--							if(index <4096)then
--								color <= X"0000"; -- RGB : 5-6-5 -> 16 Bits
--							elsif(index >  4097 and index < 8192)then
--								color <= X"F800"; -- RGB : 5-6-5 -> 16 Bits
--							elsif(index >  8193 and index < 12288)then    
--								color <= X"07E0"; -- RGB : 5-6-5 -> 16 Bits
--							elsif(index > 12289 and index < 16384)then    
--								color <= X"001F"; -- RGB : 5-6-5 -> 16 Bits
--							elsif(index > 16385)then    
--								color <= X"FFE0"; -- RGB : 5-6-5 -> 16 Bits
--							end if;
							ns <= s15; -- Outer Loop
						else
							ns <= s22; -- /!\
						end if;
					----------------------------------------------------------------
					-- (5) Execution NOP Code
					----------------------------------------------------------------
					when s19 => 
						dc   <= '0'; -- Command
						scl  <= '0';
						sda  <= '0';
						cnt2 :=  8;       
						ns   <= s20;
					when s20 => -- Inner Loop
						scl <= '0';
						sda <= '0';
						ns  <= s21;
					when s21 =>
						scl <= '1'; -- Positive-Edge Trigger
						if(cnt2 > 1)then 
							cnt2 := cnt2 - 1;
							ns   <= s20; -- Inner Loop
						else
							cnt2 := 8;   
							ns   <= s22;
						end if; 
					when s22 => -- /!\
						scl <= '0'; -- Idled State
						sda <= '0';
						ns  <= s23;
					when s23 =>
						cs  <= '1'; -- Rising-Edge Trigger : Stop Sequence
						dc  <= '0'; -- Command
						ns  <= s24; 
					----------------------------------------------------------------
					-- (6) RGB TFT LCD Initializations Ending
					----------------------------------------------------------------
					when others => 
						rst_tft    <= '1';  -- Reset Disable
						bf_out     <= '0';  -- 0: Ready , 1 : Busy
						flag_init  <= "00"; -- initial sequences done !!
						flag_start <= '0'; 
						ns  	   <= s0;
				end case;
			------------------------------------------------------------------------
			-- 3. Check Start Pulse from Top-Entity
			------------------------------------------------------------------------
			elsif(flag_init = "00" and flag_start = '0' and start_p = '1')then -- 20nS
				flag_start <= '1';
				bf_out     <= '1'; -- 0 : Ready , 1 : Busy
				rst_tft    <= '1'; -- Reset Disable
				cs         <= '1'; -- CS    Disable
				dc         <= '0'; -- Command
				scl        <= '0'; -- Idled State
				sda        <= '0';                  
				bcd        <= data_in;  -- Latch Digit Encode Number
				col_x1     <= conv_std_logic_vector(col_addr , 8);
				row_y1     <= conv_std_logic_vector(row_addr , 8);
				col_r_8    <= (col_range + 7) / 8; -- Ceiling (ceil(col_r/8)) -- !!!
				col_r      <= col_range; -- Latch
				row_r      <= row_range; -- Latch
				col_x2     <= conv_std_logic_vector((col_addr + col_range) , 8);
				row_y2     <= conv_std_logic_vector((row_addr + row_range) , 8);
--              index_t    <= ((col_range * row_range) / 8);
				ns  	   <= s0;
			------------------------------------------------------------------------
			-- 4. RGB TFT LCD Normally Display	
			------------------------------------------------------------------------
			elsif(flag_start = '1' and tft_lcd_p = '1')then -- 100nS (10MHz)
				case ps is -- 100nS
					----------------------------------------------------------------
					-- (1) Setting Column's Address and Row's Address
					----------------------------------------------------------------
					when s0 =>
						cmd_RAM1(1) <= X"00";              -- Latch XS = 0x0002
						cmd_RAM1(2) <= col_x1 + X"02";     -- Latch
						cmd_RAM1(3) <= X"00";              -- Latch XE = 0x0081
						cmd_RAM1(4) <= col_x2 + X"02" - 1; -- Latch
						------------------------------------------------------------
						cmd_RAM1(6) <= X"00";              -- Latch YS = 0x0001
						cmd_RAM1(7) <= row_y1 + X"01";     -- Latch
						cmd_RAM1(8) <= X"00";              -- Latch YE = 0x00A0
						cmd_RAM1(9) <= row_y2 + X"01" - 1; -- Latch
						------------------------------------------------------------
						index    := 0;
						cs       <= '1'; -- CS Disable               
						ns       <= s1;
					when s1 => -- Outer Loop
						code <= cmd_RAM1(index); -- CASET
						dc   <= DC_RAM1(index);  -- Command
						scl  <= '0';
						sda  <= '0';
						cnt2 := 8;       
						ns   <= s2;
					when s2 => -- Inner Loop
						cs   <= '0'; -- CS Falling-Edge Trigger : Start Sequence
						scl  <= '0';
						if(code(cnt2 - 1) = '0')then -- MSB First Tx
							sda <= '0';
						else
							sda <= '1';
						end if;
						ns <= s3;
					when s3 =>
						scl <= '1'; -- Positive-Edge Trigger
						if(cnt2 > 1)then 
							cnt2 := cnt2 - 1;
							ns   <= s2; -- Return to Inner Loop
						else 
							ns   <= s4;
						end if; 
					when s4 =>
						scl <= '0'; -- Idled State
						sda <= '0';
						if(index < 10)then -- 10 : RAMWR (....) , cs = 0
							index := index + 1;
							ns    <= s1; -- Return to Outer Loop
						else
							cs   <= '0'; -- CS Enable
							dc   <= '1'; -- Data
							ns   <= s5;
						end if;
					----------------------------------------------------------------
					-- (2) Write Font's Data to RGB TFT LCD's Graphic RAM
					----------------------------------------------------------------
					when s5 =>
						index := 0;
						cnt0  := 0;
						scl   <= '0';
						sda   <= '0';
						ns    <= s6;
					when s6 => -- Loop-1 : column (all the rows)
						cnt1  := 0;
						cnt_r := 0;
						ns    <= s7;
					when s7 => -- Loop-2 : Font's Byte Data (one row)
						if(font_sel = 0)then           -- Full Screen
							code <= Font160(index);    -- Font Size = 160 x 128
						elsif(font_sel = 1)then
							code <= Font53(bcd,index); -- Font Size = 53 x 32
						elsif(font_sel = 2)then
							code <= Font26(bcd,index); -- Font Size = 26 x 16
						elsif(font_sel = 3)then
							code <= Font16(bcd,index); -- Font Size = 16 x 12 (Padding to 16 x 16)
						elsif(font_sel = 4)then
							code <= Font32(bcd,index); -- Font Size = 32 x 16
						elsif(font_sel = 5)then
							code <= Font16_1(bcd,index); -- Font Size = 16 x 16
						elsif(font_sel = 6)then
							code <= Font128_2(bcd,index); -- 111 ?
						elsif(font_sel = 7)then
							code <= Font16_2(bcd , index); -- Multi-Characters
						elsif(font_sel = 8)then
							code <= Font32_2(bcd , index); -- Inverted Triangle or Square Shape
						end if;
						dc   <= '1'; -- Data
						scl  <= '0';
						sda  <= '0';
						cnt2 := 8;
						ns   <= s8;
					when s8 => -- Loop-3 : Set Font's Color Data
						if(code(cnt2 - 1) = '0')then -- 1 Pixel
							color <= color_bkgd; -- Background Color
						else
							color <= color_word; -- Word color
						end if;
						cnt3 := 16;
						ns   <= s9;
					when s9 => -- Loop-4 : Set Pixel Data
						scl <= '0';
						if(color(cnt3 - 1) = '0')then 
							sda <= '0';
						else
							sda <= '1';
						end if;
						ns  <= s10;
					----------------------------------------------------------------
					when s10 => 
						scl <= '1'; -- Positive-Edge Trigger
						if(cnt3 > 1)then 
							cnt3 := cnt3 - 1;
							ns   <= s9; -- Return to Loop-4
						else
							ns   <= s11;
						end if;
					when s11 =>
						scl <= '0';
						sda <= '0';
						if(cnt_r < (col_r - 1))then
							cnt_r := cnt_r + 1;
							if(cnt2 > 1)then
								cnt2 := cnt2 - 1;
								ns   <= s8; -- Return to Loop-3
							else
								ns <= s12;
							end if;
						else
							ns <= s12;
						end if;
					----------------------------------------------------------------
					when s12 => 
						scl <= '0';
						sda <= '0';
						index := index + 1;
						if(cnt1 < (col_r_8 - 1))then
							cnt1 := cnt1 + 1;
							ns    <= s7; -- Return to Loop-2
						else
							ns <= s13;
						end if;
					when s13 => 
						if(cnt0 < (row_r - 1))then
							cnt0 := cnt0 + 1;
							ns    <= s6; -- Return to Loop-1
						else
							ns <= s17; -- /!\
						end if;
					----------------------------------------------------------------
					-- (3) Execution NOP Code
					----------------------------------------------------------------
					when s14 => 
						dc   <= '0'; -- Command
						scl  <= '0';
						sda  <= '0';
						cnt2 := 8;       
						ns   <= s15;
					when s15 => -- Inner Loop
						scl  <= '0';
						sda  <= '0';
						ns <= s16;
					when s16 =>
						scl <= '1'; -- Positive-Edge Trigger
						if(cnt2 > 1)then 
							cnt2 := cnt2 - 1;
							ns   <= s15; -- Inner Loop
						else
							ns <= s17;
						end if;
					when s17 => -- /!\
						scl <= '0'; -- Idled State
						sda <= '0';
						ns  <= s18;
					when s18 =>
						cs  <= '1'; -- Rising-Edge Trigger : Stop Sequence
						dc  <= '0'; -- Command                         
						ns  <= s19;   
					----------------------------------------------------------------
					-- (4) End
					----------------------------------------------------------------
					when others =>
						rst_tft    <= '1'; -- Reset Disable
						cs         <= '1'; -- CS    Disable
						dc         <= '0'; -- Command
						scl 	   <= '0'; -- Idled State
						sda 	   <= '0'; 
						bf_out     <= '0'; -- 0: Ready , 1 : Busy
						flag_start <= '0';
						ns  	   <= s0;
					----------------------------------------------------------------
				end case;
			end if;
		end if;
	end process;
------------------------------------------------------------------------------------
	color_bkgd <=	X"F800"   when (rgb_code = 0)else -- Red
					X"FA20"   when (rgb_code = 1)else -- Orange
					X"FFE0"	when (rgb_code = 2)else -- Yellow
					X"0400"   when (rgb_code = 3)else -- Green
					X"001F"		when (rgb_code = 4)else -- Blue
					X"4810"		when (rgb_code = 5)else -- Indigo
					X"8010"		when (rgb_code = 6)else -- Purple
					X"0000"	when (rgb_code = 7)else -- Black
					X"FFFF"   when (rgb_code = 8)else -- White
					X"FE19"		when (rgb_code = 9)else -- Pink
					X"9772" 	when (rgb_code = 10)else -- Light Green
					X"AEDC"	when (rgb_code = 11)else -- Light BULL
					X"0011"		when (rgb_code = 12)else -- Dark Blue
					X"49C0"	when (rgb_code = 13)else -- Brown
					X"8410"		when (rgb_code = 14)else -- Gray
					X"F420"	when (rgb_code = 15)else -- Dark Yellow
					rgb_color;   -- RGB : 5-6-5 -> 16 Bits
------------------------------------------------------------------------------------
    color_word <=	X"F800"   when (word_code = 0)else -- Red
					X"FA20"   when (word_code = 1)else -- Orange
					X"FFE0"	when (word_code = 2)else -- Yellow
					X"0400"   when (word_code = 3)else -- Green
					X"001F"		when (word_code = 4)else -- Blue
					X"4810"		when (word_code = 5)else -- Indigo
					X"8010"		when (word_code = 6)else -- Purple
					X"0000"	when (word_code = 7)else -- Black
					X"FFFF"   when (word_code = 8)else -- White
					X"FE19"		when (word_code = 9)else -- Pink
					X"9772" 	when (word_code = 10)else -- Light Green
					X"AEDC"	when (word_code = 11)else -- Light BULL
					X"0011"		when (word_code = 12)else -- Dark Blue
					X"49C0"	when (word_code = 13)else -- Brown
					X"8410"		when (word_code = 14)else -- Gray
					X"F420"	when (word_code = 15)else -- Dark Yellow
					word_color;   -- RGB : 5-6-5 -> 16 Bits
------------------------------------------------------------------------------------
end block x1;
--**********************************************************************************
end beh;